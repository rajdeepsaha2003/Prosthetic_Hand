PK   �kjX��vr�  ų     cirkitFile.json�]K�۸�+)�*��$ȹe���Ʈ8�<S*�wX+K��w��@if$�Z�Ќ����F�����j��&��bV�bݘ��l��jrC�tr���>��L'�jޮ�6��~r��}N�?LR�??�Wf��))����,
��(�L-xb�LBd� ٜLn>�M_ܝ�3\wn�{;+c�,�d!T�^�D�&O�eZ)�JYϽ�,҂��JDjt�sQ$Z/�bi�x!C}�j�IH%k4�I&8I
�
JT���5<��D�<OD^�$/2�*ʒ��+3&��T�A]Z��<ѥR	�i.KY�&�/b�f�fd�N����ȠUF��B#C0�9�Bj�����(2�Q��/��C��D�I�%R�9]�$cKȂ��½�B�b]h��)jh����������bS�/$����n���!�Rd�`� ���Id�U��Z�*g�?�	]��.��t$t9�<]�����14�m/9�С�Unw���pU�-F�(�������֪"�,�ȡ�F%�4%2KL&�ݠ��.i"9-+�y�9D�BHb�'B�v�r�dDd�����2�����B�9fd��fhԅ%#s�n g��t∡C�n��ti�%��}@
&��%�v2��t�R.��U`d`R��<�]b��y&�С��[<�
c@Z�9�_�bd��O?V��A�X1�3������,"haQ�p��`Y�W-�i���+��"wQ)BK��$��E�lQ�B"�dNK�3�-y�Eo��8�<�G���p�Q���!$�\NT�q*۩q��&�Y�H18�Y�8(f2���ĈBr���ik�8j⠘�A1��b�J�A1��b~����xD�fQ�/hB�n��Z��++�#���3�0�zr��OpX`.��6L�3ah�n�#h�m�#h�l��C�`�A3Z�A�S�'h��G���	������
4�3�4/3�4�2~r��Kƣ4�11�i������ش�5ؔ��l�F/�)	�E��ED�"�hI�hQQ�dQ��qP	�q�K�����/�`�4�i�8 �qP�⠘E��qP�⠘�A1��b�,�Y�8(�qP�㠘G�qP�㠘�D18%��rr��)	����NI൜�/4%��ǖ�+NI൜����NI൜����MI൜����NI൜����NI�j�$����x��}j��{�������ʧ��uc6�.L9�W�uS�fr�	s��4s7�ܪ�:a���eԘ�`̞�R'�D6��F�U`dஈ�s�f�{arc��a�&��`rp���nh\�Yhd��։��X�%��8$�q�]/�4�{_�i�m�ѝ�>���#6����%�zU���'k�ۑ�;7:�,w�[������5�5���+Gxz9j�k���%x�9n�+p�Q^�z�A�e�x�Dt܀��x���rS e��(I�� ��� HY/7P�z�) XGauSn��S9���u�/�s�Zۺ�Vj͑5Z������G��P�#)�R��sN:T :�v��.PK.��-fG̱�DC�m�wW��R �
<F{=F7�uЃZ�AX�2,l:$ca˰�eX�v�Y(��RX�vuY(X`r,09�M���X`�`��`�\p�9��.p����.p����.@��EY��Z����8�2-����9 ���-���
.���R������9.�9���9�I ��,���,� ��l����9.	�9����"����'�Z��.t/'�l��N���g5u��%V��%L ۵{Ə�1�n]���F����炂�V���햫� u��	S'M�8u�]j����`�n׃���`�s=���\�zp׃��3���ٵ]��=��ω����N��4���� Wʠ�z�u���?	C������0�2���|����QO�B�=���R�!�E=]Y9�����
&���8Y\�0R����+��Z�[=p��Cމz���r�Q����cy�u ��!�B�!W�9䌸�Pb��c攀9;�܆ ��G1	�s���P?�>S���&���tL�*���������B�Mt���Ml���M|�$�Mb�$�Mrؔ��a��7�aS�oʆM��)4��٠��O�1��8�?v��r9_4F���n\Ue��/�M�Я�L�H�Df�F,�I9MDIS��Έ��6����lm0����TmǼ�*�r�����u_�o��ikӝ�>?��?N��M�ԫ_�'+��}v����ܺO�/��Ъ��L��6���V�z'7�^n�mܘ�c��K��]c���ci}k���Y���.�mc�1�,��������n��}���L��\�������tgf��[T�),�3��J��>���V:"w��V��]��y:Y7�].�3f�}�_uS,�~?%����2N�O�<� �ّ�MJ��`/N��8��6qy`-O��(04e䨉4�2�$(	),8����m9�R<N��a7��x�|���-�P̻H1߂y�x���Bz|���-�G̷�C1��{�| ��� �zb�Q9K!r�x���E�y��(aǂ<��'8�xׅ����C�-������N�����@��'U�L(BU��>�ϔ�lP�}Ec���2\�i,m���X�d����ʩ�Le?���v�XjEg�f��v�R�<��2{��G[�bD�X'fۙ�gꠝ(w�۟���Ws8����־h�������<����Ãn~��v�vF��H.���4�_P�1+�i����Xb7�2�ژ��)������H���;��B�8��+�'��A�^��!�����m$q��1��bJ��c(ѐ��I?�;<RT���NG�a��������Al쯼��I@?��p��L�s$鷤$��#v\ v��b�W��;����Uz-�C��LI;;�L��O�㙕�)g�[�n/�2)�����A�4)1ʒ�E�H�@?�fN�S��/�߂������%~�:����KHEYh��pDOA�
���PO]x�]�]�k�6HLl<�كt�����+��,�j��u��;T��_��wo�_rCK�:���]�8R�j�tqoʟ�R��Ӷ|������	�����I�0������;n'�[uӾ�W?�]�ˋ*:mfU��wt���CT۬¿�3�a]������t}���������k���5���'��q�k��>ϻ������B.��Rj�e�y~��Q��I�8�ᑺ�~;�nay�݋(�B,�1biT���5��l!�!;����@l ���01!�"B�E��1b�?<-gB_"E !
*�N�l ���@����@���1v�i ��aݙ;�����|��\r��=��`R�7ܥ��$�R�@�DzR��ٽ�%&�ְ2�ȰPX�a�O?:�,�l� �x_*���;�-5��L�{�OL(raE���ȡP<�:$9(v��| 
pd�K�iCw(?[
�ݻ�b2JXT��hG&��x�u��I��	so�J8}�X�w'��R�ӽ�/&4`<V0`x�uHhhY�r{��TC��ֽ�0&8`Q���>��a~r�P1X���"�{�dLp(8@7�D��n~�1�01	�C1?8vo�	��>���A�q�uXpHH��K�RX���"���Qs�0t�n���C���9t�]ϳe�k����].`7��.�0�:p�`��].`7J�.�0�:p!	���eC�kC�ڷCܼ+AY
��P��p�]��pq�yׁ��oH��P�1C�P̏��eE^�D��ح�A����)Z?��'!���]3ab<�.p���+p�a݅��	01�P��{��[���
��ؕ����7ܺ������@��{�[���.�>�,��ί��w�/�5M���ɍ[�M����)ѫ�^����sk>o�w�'��PK   ZjjX|�<�d� �� /   images/3718d1cd-d7a7-459c-8466-c70e7021b870.png��SM6������wwwwNp����ݝ@p�� �w{��y��N��0S��5U=�����eE)��   EFZ\  �����a���� ��J�j����6��DD ��8���m'iW  ���ܴ$� ދe�E�=O_�(�RE�TJ�j���(�����I.��k�����8�|0f���s	��mP"0�L?���z�=������=?Ⱦ�q\���,��� ����]\\�|A��7��KVS���U�<��u��4����*j����6��#c��Ǝ8������w�PL����ݣ���xb���Ҥ���� ��/�]ɟ�{�]�O���ș��ʛ��F�1J��W�1�L{5�9�1sURtY���7�U�q�qۓ*6H.�&�1n���"��E������|�SsV�ZG���r��y�ek�������/4��cU��>Bg�@k冰�"��3�����(&,/�(�}��^�\���0�>���Y0)�O���(ޖ��"t3�~� 
�oJx�_�]��=A���u����Z��-äx���}���a��r�}�5ۡ^�j÷5G�&�v:
@�ъ�&E�0��W;D�����ƈX�`���{�!�����L�J׃o70!8?`"�Hj��c>c^G���<��7	������D��GE8}��U��[�7��Ւܔヮ#�d�ܽ��H�]���gN8�a�t�l�e{%C���D��(�f띹���	����n�P�W(�Q8������A���1������.M�8j�+:�����c�%��r}���}t��;4�Ҁ/�����䀸8�#�q��2&�4=�Ϳ�;=.�sN����ʷVF$C��9\-�A����G$k�jnQ�\}���^eVA�]����k��o���^����Ɣ[Ї�ʀl(a����6辧��<�x�G�]��d�B_��� ��$y��7L��#��}-&
��fɐ��>%e��gܘ�nnN�Ah�m��0�oaQ����.���>�'�.D#�����b˧ӝ$��+J=�#"��K�ֳѥ_��3�[���ԋ8��L�$v}SkkB��?�s������2�P��U������7�g�9P`ŀ p1eL�G5"�[+ ��bKqGR-˲=�.Q>���^!7�Z��m4A\��u���"Ii�O�g�i��Ɍ7�� �$8�5R��<�Q�
�H����=L�V`�N�z}f�`R�Y�u*�@}�����lK5R��~�T�i���l��zX���S��m���
N>��zW=�#)���⨴��&�N��%�E�Q<��L��Mވr�L묒$(
e�U�SU���:��!i��*���:Y�����K���ҀJGu���
�"�O��;a�sߝCK �^�gjn+4���
H�G�Y����4r�x�����	�.h�H0}��&Q�$���F��.$�z�B��n取��Ə���v;��n_
��l*:�*Ֆ��ƍ6����w= =Ú���EJ�D�t��o~g�S�n�|�[2���J>6�cޱ�.��,��)=�MBPU���o��r�lel,����êxb�Ȟ�a4k,����Ӳ�.{w����WD�=�i"To[��5�?��@�RRR�8����-v-��j����{h�@���b��=#+e1L6v=�t�?�1�Ie��98�j�-��Ib����j���E�;�2����,wBf���5ǕǬO�cv�y�*?UQi0�MqA������C����c�g�^����f/����!]���~f<4�M�Ax(��H��a����H-��&kkk�����U<A��X	���"EA����h��ۿ��C�6<rNAX�� ?%�;6j�XH��J�x%x��<U8" �8!<7����{82f�.KN4 _��d_�6�V:=����\��}X�z�Tkw�r�%L�*,jU��e3�w��8�0�[��u�Y�E����(\�\��_�v����{�?�Q�D�SEB�m�;]YBo�:�Q�J]�T�ilʶ��QG����~�8�����n-P�<|JA�%N�p$�g�O�?\��҇���1�D��	٦��]���@,/���N���,P�dc��#lhH ��4���(0bO0�-���!�j��~����>wx?�~&06Z\�P��m���,�ص\���=3�u�+ �GCAL���dP0���FJ�K�0�p��3� �x�����E�ɰ��5 ��4�o�idG��B�i.VCaM��� �'�l(ߵ�naAcmu��F~'� 6��'����.�j���]�s��K�i�ܱ�H-b������N�a[~|1f$p�����\ 5s�l��y��'�	��NG:AR�� �A��`���7�;n��ؕ8�ԍ��6�?S�`�:���;,��&��F��[�t�/�����(���֞�J8k����+5�֬������q��i2���%s��
@ЗY4hRhZ}�6��E�t����i�h�2������WPWDD�JǗ���� t=�^�q`bg@[���.��B>��i@I��o�a��s����l˘��"O��)Ch��ք�q���	�<ۏ�,(S�{��ăψ��i�<�'���?�/�6z���-����G�2��/я唋�G�`��2�7$|�&?W�cX<gE�Fˁ�C���]q�d}R�x�N`fC�.Z�7�f��E
Ǔm���cZ������E,�OO���4�������"kWɥ*�C�[�O
������C[n?���2"#G��_�&�S��[t�:;r^���EN��$��)�Zb�qIa(,2��|�ݍ|������7�h]t��ӝUGo�up�R�H�KK�]3o��F{���'6UI'�Jя}���'�����b���鰒�i����#2��O)E�Xwpu��Z��N����B�hW@��--�a���z���5��2h(t�E�tˊ�w�/��1��h�c�e��%p�ᕐKz�c�i=�GC'iV�"�[��B�Rs�M[�|n�4�ן|�Wn���ϻZ��.-K_T`���/�j�W*��(�3l.mJ�D1a$�G�Ίn\�)!�)eRDɳԲ6���\%,_����7t|��d{��<J-NN�Ҫl���{����Z\] ���=Q/6�<1O0����~͊3���v^�Þ��w@�wJ�W��^�3v{E鞐6�:�o��o��{���QQ*�n�\�L�3�4�Vb� �k���{���K�l�<,�5�*�ɲ�a�-Fn�ʆ��OH�ۊ����I�G������T��'�;�z��pY;�05uz�e�:���Z�z��~�y頺����JV����!5�=E����ѐ�0^����6�d0�6�m���<0�����%�̈:�[X�!��4�T��܍�ҝ%;RV�"y*�l�Q-	oXR�����sx�:гfZ��/add~�{s�Y��$��`A�uwW�n��+�����vjIa=�����u�dd[�`��r1I.���­W�e�YT�Zu�;����{�T3�̞TD�$ߌ]�A�����3���������]��J����HE]ճJ	��SB���X����׭NR[����[����������;��=/

�X~���V���~HPl v��T�Gv (�lU:�ĳ�v������F��+i�1e{s�	KjGKb|�2IH��yr�|�~�P/N'�o��������V�[����9@��l�� ��{|3���E}�s��ea�tu뛛��������~]���jP�,���:�w��j�{�# nj���l�]��7��3�y
�fy5��t��ꦜe��4c�?!�4��zE��%�d�5�{�G��ء*G�"P�bW��L!^�qn�Z�\oXg?^E�_L�4��	]#�@\��>�	�+3ˆ�?Ε(�Iݕ3@(P�W>�0)H,�uF+��c2^!��]&zf���:-�'������!U�I��6���nN�6�?�5S`����L���\,���-VʌR�5��V��Ơ��B�E����ɿ�7��,۷럐J�vȻ\ 6�L�����ŻWÃ<B�o�Z�(Gw�q������?�pĉ�i��Q-
T|�@�L��#"^	��;_k=���Ҭ�:�j��<�����݋�ِ���<�����C�]���Kqo�*~8���<e�!��ѭ�p�:��	��[���#hH$d�����ζݫ�~]T�g/���� ��������-L�0���Q'�Ce� biG5�T��B]ŗ������嫅�,�x�>~r�S.�^�p=��п��DMeC��w-6y�>�G�1C�K��(�I�3���FL\ Ձ��r�^n@���dO�tm'�F������'֐���==#u;�4 ���X��m6�gEϿ�����H�߽�/AH޾�&Pi�Z���z1z��y�)?#&]kWx��j��:��n�-4�Yt��"�ܻW�H*���7����<$�st��rJ� Q*�D3<��,،(h�k� �?��ܭ'A�AFd�h?��`���f�o3.�s�~��IJ��^0 Za>I,x�L�Mu�n��y�W����8��x���#�JzX����o�Ǖ0����ī���K~�|�Ib������ uC�~G�#e.+���뜃}0����]�ȴ��E�/���:I}r-�2PS,4l�ln��u�ԄqC1x_)������(�L��7���Or�U:9m�����j�*��X�N�.ߺ_��އޢ�O�m�z���Ϥ�W�]�IWf�;b�%NFG<70"��;D�����q�^��tȬ� Y_mv�'n7�;��<��B(���R�`P⛡{6|��!��zj|�'��`S��E�%�&@�-��ɟ��2)��^�vA�ß��u%L2M�E�c_V���h��6�\�(u�g,���:��sI�0��(�r@����f'��M	��P/������
#��)#�r9����Qж���4�(߳oB�h�D֤:9!�f}���P%xHR�?T�a����
�S���}�Vs��~Y�χ/�b�$hտ�h�\��RS������n������R�֠���E��V(����8,��F�g��٦ᒔJd�_�.K��AG㎷g�ݗ��F���߁zH`���9$\(�~�j��	P0%������؝�U�c�ݿqA�q~�n ��Y�����Y���^��D����)'�U���2�92¹���6��b��/l3ŝ����D�|G��N��F�fY$&sMH��j�,$� �Xz�J�D��{*�>x��qU�tm�J���]���*��̫����e������?�V���u��]�7�٭���08'_�9�wM���8���B��g�5Վ�O�v�\�<05�G����l��6T�C"
���e�n���Ӂ�U�#<,���WR��:X�a�n�Y�xz����-�KY�����0�і�&�����Ym9	�,��pV���2��T��4�y��`��"�`/�A���h�R?. }��� ����S"�����'+�^h�}��ӄ}�{����7"������H�㗣e��;G�<��
��e�I�ܷ�ԅ�f��t�Q�ohx��#����귋p�Z��X���*�n����)7�����B��34�{t�?.T�qў��J�����
���PP}=��g��3h��
�躴�̒�  0�KS��9F�ZJ|R4X�-5�H�{)I�-���F���������+���S�Ls�s�9��8���U�h>x����������t����HN^Nkai*��=�}�C6��f��3�4O^ ������abڨe��M2m�DƊ���+��ND�M��r��*�/wex�}�vt��B�$��m�]H���heB-���dZ��$| ���o��c��;�D�����`;vws3���:��1�@dĵFR�Vd�ӂ��c�m���V2��?ʪH��8S�X�6�l:���j?7%W��Eߊ�0Q+��@`M�/k"y��E�n�8,r�����I��3�F�qX�м����bD܄���qx��]��%O����.�_�t�k(���l�J�W)e��0"����+Z��2>g�L�?�0P�N�D�ojL��dV���9���{j��Q�c�<��� b�=�7~�xmDr��W��dr�@�ʗ�7��x88/����r~SQ,��1쒾���i����Ͳ������i�R�^�K��?��y��;������<G��߂�*�?K�-na*Fk�&w��<�֮.%B��>���� �]6����*���o9���R�&�qQz�z�`���wX�?k�Ү?Ƌ$�
�pp{^�A��1g-��z�J&J��Uv��|a��Ggǁ�;�*��(v��.�x�f�
4T�r�f����!u��H�g�)i���\^�P�e+�2�7.I���tnZ��^uh�KwE��4}+C+ߑPԙ֫'l'�YZ;в��đ��*�{U��ל<A�|n>�T/53��'֣oS4!�o��L~O[9�>F�xÛ�Z�GPengW��]o�'�����uq�W���äc\z:�bo�NဿR'�_:y���H:�[!�!�<�����nl�
�pg��v#e���ܷ��+W$tAJ�|�E�nr�B���+��ٚ� ��`{�g��FS�������H�vi�-�)��* q�-_(��"
>_��[�\� O'�z�}T�#����l�˜�{�Yv��J*O-�J�KɀeM0�4���[�{��̓�����Q@����s~��?$t�:�<6�=�Lf$�d�;���seWpw��$�=�Dz�*Gf�FE��D�fiG�۵��f�M\	{��2�*]�S9�k���ρ�A�Ԧ%%ׯ"K�| ���Sg�ߦ&ק�Z��Jw����XɂI/�"����m��+4�p�kl��%��}�fu���ԮNu�_��S	9ù�`���YX2?�-�mR��ol���p�d���6M�4��[a��>Qe���T�|=i�]g�{�����9_����@䞹�M��>S���H�"��8���B�1�u��%�l�dRr|�e�+�'������rE��TJ��o $��<>囯�碠� s��IP��^a�B2�-/�������� ��F���C�R�������0�7$��{N��E�g��|��Z�cyi:��XMH�K  RW��V թ��4D$S�zZ�,������MX&����h/���;p�6�o���H��ʁ�<i�?����
�9B��� ���E#+�n<�+͞��h�Cf�i:6z��
�zY�̌���> {;p���F X�{��78�F��,��]��<�Zºp�l�D�I��l���;��3��[�Q)���턇�>��uD�d�޾��.}n������W{u->�#�YFt���1�q����8�己|^BO��E�mf+ӣ&A���xm��+�an��(\�1
�C [�H���-�Ii�@�h��ِ��  ��1���$���l�\[X8(]]}��?�Sڢ9��W��#P�IQ�&Q9S��]�l�-_�;����*��[[�Bo
��tp0PޏT���I�Q)��"��U)Ə4���\���[b�����{�k���KB^�9D֦�="�˗��0( ��Ȳ�f,�� +s�D��ϖ�4+#_�;�T�_�>)�f:s�y}��ȼ�B��V)B����.�; �E;Q�z۟˗����XՍ�q���OM'MR�NB7m]��~)�=nC�N�=
�Ik�i(x�?$���Q�jxh�l4���!bWr�0,0ܘd��YU��9�U	mv�+SQ ��*'_����,���i�5IbO�Gj�G���n�_y��K�}��姱�.�J��1V���aM��z����704�?	�H;� $"Y)��nY�����=�ǩ��[_�<sm��� Θ�ø9��H�ؾ�$�WǊZ�|¦=C΄����G��&aF�X���6x�m�fx��on�ؘ(�\�b�C���E=y�֠��Tz�uY���q^��Q�!����FCXWl 4*�لY#��N�WK�"m/^�$���Y���㾌W��Ũ���Γ��Ǥ��)��2��D�W�i�	�Y��q���Rh�[�hFM����K�~jp��-��)z��6��w��]�wЗvTÔ0Ȭ�?��� )X݇�o8]t�L^ӡPݤ�F���\8��mH?����j͉ `���*|%���K�GA��F�rm��=ʅ~��V/߻7ɤ4UR3W���C��S7�O�N�,�F�9:W����h���	���V�8%:�4�rb]5ok�+��]{��ǎ�|>d��0�1R���A��@�͹�����x�i�EJ����r.���]��፳ѓ +�ُ�{��0W�̧�����<�J �G� �'?�z{z���5}�I��4������W����y,h�6W�l$�(�!#]gZ.�S�V���Q/Q콁���� ����D�h!�8�o��4�$>.��W�/*>y�{��.���s��C �Y�<�� �C�J��Z#PN� ���n�0~���BƑEw=Mw��=@���-q�J�J�n�軠X�)�Ro9���D��~���(39�ݎ�LK�5m�|���>��ɀ�;�� ��cE2�cA�����k��OB$��Wг���Ν��Š���I��S�6�@5ɲN��8�+�O�V9���z:�v���&���k��r��F��{�U��O����Q[��=k��_;I2&(8�Y�V_��}}��H�[}���w^��f�b]?A��a����I���0����+��EK��P��k�/e��dN���	�	�ޅP&���,_�����>��p{ ��Ć#�t"c F�����^��P��q.�/���Cq4oX����fH����]�}2/����'�G�b#]!õ��$��)#`���3!�Q��D�&��ܔg(¿��<X�~w_��J��tBJ���a�Y�Y���`t<"���ub�������o��1��U�����l��KDP�A�[�Å�^����؈�y%i.r���$�\g�aZ�XX��f���+���~�7Y����X�mL���x���疯b�!Tf�6�| �[�5�:v�,�(���0�"����ݮ4Z	�@��*�S|����8��#:�/��<d= �̾�����_���I�Z�`h2_`?���-)�1����:�Ѩ�K*�U_�v?�5���wpv��.�⏂�zG45 ��md8s�2��2/Ft�Is:���n��h1M�ׇh���SV���X��XpL؍+���0��-��6�߶��EC�ʭ�vFdmQ��Y5�a���c
�R�s[s������L�[R4�b���z5����Ӫ�:l�lx3ε$ĤI�?{��|u���&r�OO(�>&>�/¢���pc�0*��;�>�B�XK����(�	q��/	h��m̶U�Ϝ�+�k��>���xx���+�"s2PJ�XcUJGl�z���&԰?(7� �1?�;���Y���}���":�:�r���k��1��� $I�&$I
�t�Z����v`�Y������(������<E*�/�  �/�����%�p�\�{�@��>B+rO	/j�.�T������n�.L�a���&�]~�f���R�[ ��y����Q��P����"{$f�?�ڧ1K7;�0:6�������KBS^��������~���)�[*}���t�|7�q#�41�:�RǄ��R���`+��Fë���ɛC�N�Ɲ��c�{\����m�u��$�d����������A�`�����Ms�?��-�m&��K\�H���*Dv�n�{X���Ӑ�֮���ۦ��tk�ԴRv��^���j3gk�l�A���5�����e�fE.p(��Ԁ�բ9F�܆�����jxoOlۆgj�SqijM7-�_�����t+�O�?ޝ�.���t/o��%�������#l0mXBB���B���JL�a�Y��zP%�u��ǳJ���̿�&�w�c����є!�[Ah�+qB�9{��J:���[��G�|���9s��L���S#6�f�c�?�4,�2��-1&�Es�H���La�@9�ܰ��$4��tTQ,�����;r������V'%�#-�@�V�A;��)G]ç�V�$�j�F���"u���]�&��ΰI��A`����m�B*n��BH5��������Ĺ���_��K_$�D��c�ES�}��qÉt����!j5g7���ͥ_��\T�M�nd6��u3#`��c���.4�Y����k�]L@ћ�
`�8��=NGy�K��m�Z��{������y1x�6R��6v�-�+]���_?����
#�fp�|��vV4�����=�+T�t}'�|?��iQ�?}n����Ό6"�G�93yT����Q�$'E��E�k�2�݂��&	��Y0�X�8��3eQ�~��fp�@M@#A��W�f��!X[��G�a���>�F#��92k&U��ݍ���z�$O	jc_�L,U�$�A/,�_��ck�@���F��A��Y-?�8Nw�m���=��Ug#|k}�^��K/I{z�����#��<��%�|�Q���$.TS]��ꬊ�v�i�$�C7Y��H��ww��<B�yǕ2W��a��2&�ǭ>k��
Y-�fʻaӻ�+IY��"蛊+f(�&&7t�>��	���9�B�%��uR�����(Չi�F��	���\�'�#�gBl�:��{�^�=��o.��+5#5kR����}1s}@LY����WxY�U)e�g��
�~�7��Gh���:~�QQC����̫�5������hsz����W)�8#��Ѽ��̿�i�oW�)s.�@���8��b�����0a��Gk�D;����3)(���N�-�m��#r�?/갂��F-�b4!©9S~a�`�d�B��A����j���a1x<����SjRq}��l=�����l�6i_HM�0\�����Y,#��@H ���3tɔ���w�+�?�;W��R0�j�;!¾��D����plv�2p��nC���%ϔ��]�2ǹZLp|^�z�N��JnC�_d#6��^DYp����*�H?o�i��.̉���Ql��F��:&���\G-��ލ��\S�+�
@�Cwt�j�)��7��y���4�`ł�C����*�l	i
�s�Oq[aކ���hxEѥ5H����m�iJ-�B�u�/)~��\�Q���גx3��n�kجZ�9(Ѝ�DÜ��j�f�h���BCOϠ�̕pqAlj�Ol���&&<!����B&!���2N�][�}72����Z)����`�����V�_�����fhծnE3+�����;!�ʂPH�;j���OT���ߗw]|w���T�1ɒ���`�0M1�1�!�3�G6.��WҐ���Q�;RIp~=��x����+>)���:�D�^��x��v-��2!7#mg���E�^�QSC� ˹�!ŀ�ź�R��*)H�D�ϲ�K��7�07�	tZ�k�;Z��ɡV�����]D�,Q��R��:�}�r48���qVU+�BՇr��T_}��$Vv�w�6���¬�5*ehҍ#gh��7W��!Vʝ�ٝ�<��b �܁U��e�ʥ]G�����j{�oT���fgj�ȍ5p��c�9���U����^ ��R�2`ThX�ͦ?��t�\���wl/��(i����lT{4ۙ�3�#He��"������ ]W����Z��{`s,�C>/��N�bպ6�����l�:A��å�Z��8ꟍV�����К��W�E�y*jF�G�*v=���Gw;{Ǖ�=�U�*�#}�ar��**j�J�sV�:=w��lȋs^y�
��#V�����4�=u-�MlwM�,i��{3�*.O����qL��J�S��%����iU2��3�Q�:�<�M+�������_WvPX�R@��6�$���� -E��UVv����h���FU��$�Oˎ$�����+�����e/����+�ٰ:���J��^��q�Y.�e���|�v�X��	�s���]���0uHl�1���<YQ�+��9������5�x�Q}f�R;Z�blX�k����ػ�8'he*ﲲn�����kw4f��e���}��Z걂����:K`�'h�cq�M���������ث`���\7W?��pu_d�8?��u�[i���&+��"�.��hck]�� J��&� ��&-ʠ��\�ݛ�B ���%�%]�⩭�C���lmT XW��f ;Ac-ś�N(��\�d]�8��9}�b`�$�:/iK=��%��wxi�p1�:�1�i�M��fU�ˡ�x������Gb��iNh�4��d�����\����={�����}���R0��T���4m�{��- �|윪/�O�D$�g|�g+S��+�rߪL$�`gB$�hy_���h+�J	9n��лx!�y����l���R,�	�����g�9��	�t��,�-R-������ćY:c�D6$G[]�����8���W�7�7"o~`�4󹸨x�q��|��~=��y�~,C�x����$B��/�u����Jg�Zz5�����m	H��ov�fdn��:��UQiD*�S�G�`̴-�>����Ĭ�0$ĳ��� U9�+��\�$�:�~���/06Ʋ_35�/�]���6&��u2�oii�����Q��18�nl��nۜv��ԭ�h؁�@ ,T�GҜ�Y2��c ��}ވ�hh^�/hZ�<E|�G/<^B�4�*�B�D�/����z�}�G�%�����9+��oy��ޝ�軹�R���7��B��*j��fHǪ���/�]Ug�1�rFlP�}�_�I�Vg��¤�e;����XR��RN3�rŬ��lx��7�Ur s�r �,�K�8��V�#��4�_�?d�'���w�m�Au��0_�YB���ElW�O���n��C�J:��Y|31�+l�� f�Cg��3�j�*�H���}ӄ��	��qZ���`�\�@��9h�~��h����ս��ٳwwA�wA0��U�����\R��8�ߜ�nJJՍ��C���U���	Ȯ�fb�1�}C��SQ1�)Z��� ���uu�9}x��t� pN-R� �X�6S�#��LtH,�JL�]�� vwZ�:�G� 7���
�L��E��HBJx�n�y�����Q-L��o~��8[����xx��=�#�99��6ڜ'ɰ��cX��9��=�+�J��\�w_c�@�1�(��8�wF�_%�o�X�%O0~��PY��Ň��v<2�&��Jvͫ���"� �����P"3�n��:6���ζ$�����{�Ѻ����zK$����S�iu��Dj�a�s3���)�r��֫���N[<��0�(G�b�YT�;�7e\=I0�8HI���Q��fpl��;<�Ǔ��OaR��h
������b�P�à;��)��;)Z���7���eP��n>m�6�Q폧�;�/էd�*��3��&K��=�#��J�N���C��}ǽ-�L�X�}+`��.O�T��6�N,�~l�E�X�f/냂RKt�h#2�l���-�[��@�hϻ( ��k}������� E��B��d?ݶr���l��,�=�B|z���^�S=N�!�S���B|t$XO�Z���6R�7)�r�J/�۟YZm�����h�R~��6���u�$K�!JM��MO
K�^�K����o�5����Ѵ<���Y1���q�V�-hn�*&�!C-�Eqb��9+�6�!�Jώ�^B���Ş8p��!Br�@�P��ƭ�A˂끃�q���x}x��q�C��%i6���ѼѳY�s
��<�5}@3��Oլ������ĝL�}Yl��T*�jW�����ea� }�Y�^���y�C�c��Xd3��Fw��_oR���+5�"�g z�7���2 ��o��8����y|�;�Uj�L��aՅ��>�x�C�G���:55��ae���]��HzM�������?���GE�r,��������F��?u��'uc��8���E��^�/�T3�=�	��II�v���:�Ϩ����T���X�
�d����~��y���r�/�He%]e3�.�O7��C��JW���)T�,��B9�n"�<]
�{LH���`#γ�f����tD#��}s7��;K��4���V�U\��k!�txMU�JX������*Sy�Ѫ�����Y#�����[�RGW/)��x�6PԆY�J'��:g�<y�������+���@���Owŷ����70�����{ܖ[sgc�P�:<Gq��a�������/)�7�'�g+Ґ�����Bus�JuWhTP�̚�;z���f�N�fkuC���5��D�ռ�egc��93� ���t�pojϯ3�A]�@��ݰ���'�ooH�c�n?]�'��z��R��z��4��NI�j��Q��'����O����ؤ�ʃ��Wnt�{��"!-M0x��T>Z8�k�>J<��S����3�ܜ���D^RoX��x�x��a��ܫ�6�:�S��/� �2;$���SSH�O��ŭ���
��v����r�=���o#؅Y_�OW�@�y~�w���<o&�������p�1����cP���2�$���A4��B��X.��|���c
]��[)�Y�Ox�=d2�@i!<ܓ����TI�w�U0-�'δ�iѯf��j�#) ��8�|�9q�5�|��Q�6^~uj���#��3���v�`}q3c%GZU�H���L�F>�ڡ�����A�X��J/�]�_��q?b�Ah��ݵ9`T�3���Y�i���Q�H,k�������'���=�����l�m@oO��n�c���\�4���nl�`;j�W�dv�5Wѥ2=6YQ��P)�y��RC<���p���M�U��,�����+�%	��P�@��2�_�y���Ef��>�U<��Ymq�v6Tuj�H9�h���Y��y��\��t*~}V�3��3u��ʩ��^{���b˹���4q^���ZrعW2qo��虯������;?V8��Mu��G��.�;d�\�p��"�''�%a��=7�u1��ۥD�?F��$���)���%恹���\���B�>D�D��y��oۢ�.��Cl�Rc�W	+Q~a�)T���jF���7���/�V��*J�0d�Us%�JC(�����j�������N������0?	Q���x�N|D./W�&p��YY�Z�E#Y�>i[j)�%(t�0��a	��d���?�D'k�r�t�ݑb���{���׬�e(�d��b6�)''X�i�تm���5��TG7�����A�a�D���E.p�(RO d ��G3>�Ƃ�j�&Buo����=/��%�\[��8�a�Z��S+�rH�����:
/��y\|^��	�RRVΐ%����P��NjH�T�*���^�
w�BQ6��mNTH����1}�oY��NeE�J��4��w	�k���a�wĬ����#	v2�u�'��M0W����
3ު���0#���*��jͧ<��H�|��y_�p�4|տ_�Z��7�!W��Y!�Cv=c�q��j�f���c��i��wu�ڬ���%!�.���bP���>��/>:��+�d�&����&bɁ�
�A|J�p��ɠz��U�YĿA�ҿ�13�V�I]>��S9|�**R��s~"�8%�ɡgT�Vl4 6|�]�-��������9���\��~Q�g*�Z�y��٤�/���4���#R��XԆl�\8x|���}������S�)���pS=�C�3q�ea��T`4��Aӂ�}ޯ������[�*��B�䛫rn��n�9���W�
�s���^*�ÚKRnT�|>��T Ô��]��{���rs��i��P�@�x�+Imo��/|	)&Nl�knѮ�rM��d��v���x���wh�����n����/��/�/��VV�w�j�cZ7��鹪�|_u$�e\.����5.�EA7�nz2���xuvJjV������í��a.�pڟ�i�o�2IK�n� ����m��P���E�oe}��Y;ɫS�[�5�>����v�&���_� ��1�	!��f�����Ur-�ͧ����U_<�_���w�Lk�'�hVV$��?=2����T=�y�z������I���_��N5`�3E�#~�%�tLq0��b��+6�'�rwq�!ݢ���|��,�a���}� ~@���9��B9����~���=z�ȟ`�xKE�qWO`�dէ2�§QX��t!�y/-4�)�'�q �;E�Κ?m��m�b��%�E+,,[�ϵ 	����O��Sב���g{2 ?F�4��8��d�:�ħ�"�G#@����%J�I�iu�Kwl��~�����𫯭4�Z�Q�����`Ŋ`ڨhվ�q�h�BϺ����(
TOm�/�" [�QG�}0���-kllȠ|U��F(bt1��'"?a���!��Px�8��Ϥ'������H�P��J�"J��#bÁ���l�x�G�����[�pɊ[�fr��s6��$�>�:|��Z;��U]�غjs�����[�*j� 2�%��&K��N[V��|��J��b͆ͪ�Z�xؿ���D[Ao�H��/�#�e�!�(Nz!�ߊT��3����)���<^ouV����O^j��_S���MN�m�VV� ���sf%>�uvd�X
�>�:��Z�N�{���-���b �}�B�b�����M	��M��X�O� 9ތ4@���Q; ��7����A<����7}g$l}}�ӥ4��D>��Mz�R|N9�]P�r����� �Pf[�牜�����`�硞�?��s;8:��:�"F}ܷQ��O�E�n�T���ӏ#F�~�ꥆ����lZM���X���KW}ܑa�aN��κ>"Ƈ��u��5�/�IB�Wf��d*���7�e�S��A�ۈȒUiJt�,�O	<�؈��(�7��/�A4���pO��Q�.�?So��x`��l狿�ݯ���ݲ�uaBK�geeӁ�VAϟ��Ͽ�.�l�.���ӵ޳];��M��֐� �$�����^8oխ����I'fӲ��lC�͞�a}�.��4 F�$�t;���#�Es>:� "t� E����Ȋ��z��C��c�Ol<��O�ֽ���=���S��J��*�.���Դʩ���yjG_~m�gOt]ؾ���uR�J��jW ޑ���'Þ_�no�o
�//z F=>�T��J�a#��v]HN�ơF���m�#��FH�m��\{U�8��hr]��������1�u>M�7! [�J�޴:Sӕ���-�g�F��5�U�;��lW���Uz\W�N�ZL�?a��3k�%�E���[�4����V�\��B�W��H�,"�Oj+��f�7ң��R�-Z�Ӷ/v��|�~��H��C��=% 7T��W�%}��oC9������0"���ٿ��dy;��;O�<�[�n��BnL�(G}��/-��];`������޲%��ZSxɿs�>o��b\���Ҳ-�y�ܦU�2��	c��a��LzW����n+�.: ��0�,Vf������ ���~�ȳ�����y��](�\A��Pd|ȇ����[~��W���|���O�1j�
@ܱ'�+
@,1-Ĉ���`��_h�Xh�H����m{��a>��|��D��-`ztb=����v,#wƧ�je�d:�����eKҧ���d�$��+����п"����ׂ�J`졒E���&"<M]�>��1��D�=�(�����Ni��� �Y\��#F�ؒ��e�� �k�F���/�yx��-�������d^^]���-k2+ ��w���Y�4���S�N�ו�қ�F����$�l�j�J�V��Hӑ�<( (q�,�}��3�y�H.K� Fb�Җ�M�<���� �����@mc��������G���>c#`֖Qm�,5�ŧ��5*�֌��M'��ꕋּr���W'=T1%����@"��4]60�t�PAT	y]~�2$+�h0BJ�g��ڵ��Ƣ�x�K�+U��́��r�m(a9�^�:S�X��a���u;v��={,F�̷Y�̨�2��S�GO �ٓ�>��G�}�lIƭԨ�+��}����,����o���-c���S����M�M��u�u[�|�*����m�T/��Y`}�*�0O��w�a=�1u�Z<�q"±Cԕ�"U`E�r~))9�!���h둾�gG�ܶ��5{�ƂU����ի�[V�����ٯmG�n��ޡ�5ʚ���];�5�{�H:�Z�Y�NMr1E�hڂ��{����YM�\/���/��IHu@��q%7z��� :,�MP'����XF3]997%�sF��O9)d�<�0�;�����X:�;6�Ko�Ӗ���|Q��v����O�z�[�Q�%��$-.-ZM�x;��ȩ�����%�Υ� ~OU�ha����t^@dmC�I_j���uCVe�KI�B:(`�:G��y"��L�E�tCΌ4����O�E[���	�T�5j��$�Ϻ>j�ْ@MYa 6V�7ê�x#�e*���l=��5�=�r᢭\�fՅe D�g�L�3�0U
M%W~⩗���z��с����k]gӓ/�g���e�ߥ�D�v�SN�M9����R�����Q�8���N���/�s%�.�4�EZ�����"k>�����~���vv����ˀ4|�M�� U�D�D�-��p��y߳�e���5k;�?��g/l�z�Q�Q��Uk\ ��w �<F60�|�Z��;⿫��<�����莏������pÀK$��vˬ��!�/��4{�����(<~n{a�fե�./",/��7l�7m��9+VJ�C��;��+��I7'-��:��ߏ�P{�K�L�g�v`Ê�uYm.Y�?��'����|�t�V��� ��X��%����k$2�'4ՋP	�x6����G� �Q_�#D0���/X�߃q�Hx2"��1]avl�:>6����50�>�؁���.�X��:����B�< %��R_ņ��6�(��6�r㆝�ভ]�,I&ږ
��^➘��W�ќ�g�^��c�H�MF��{��=�J��,���!��XOI[�ჷ_+|�{Q:kX��&�S �*�jҠ����
�#�P7iA��@i٬��{تu�onښ�`my5@XQ��%��HJ���Ї�钫98�Q�c�d/��_��#��=���2xqN��?�߫4��)�����{Entd� �a���>��wn��UK7��T}*�;z:mu����<yb�_m�O�t�:���6�T��ڐ�Eف�5����Y��s;����޾k�Z��;f߰�Sw;�k($����b��w�C���Q
ր��|t
��vҜ���г3a�6[���`�8{�y�qH�1��˝�-^}�G�����?8�q�m�Z�j�K�.�]�\p�����޷�ə�Y����b�|{�/P0�eԦQ���"��Y[�;ҵ(�V_�Z}�i��%+���)۵�p���LV����Ӄ�L�)1��=S�A��|:f��%-?�����\u.6%��#`��h�	4ª�kY@��/1�.�����Y��|���ʆ+����e"�@']��QC�]�`�?��6>x��kk6�|���z$"��Q?�G���7�����=�H��ĿȞ�e�����k��&�|V��<�b�b��[�:g/Zsqі��wO�U��O�61��H(��L]�t����Ȼ�ݗKo\WY��n"V��U�Ր��*|��yV��((ْN��$�q���5;S� Wkj��_�o�[�Or��KeB�|>,��^�����E�,�O�i�Zy�����`mI ����0�B
Á��H�����xa��#�>�L l�ղ��[,4Y<�X��s{�����۷}�'@IYO�L��>xh���Y{wG|�T�PHO��R�6._�U6o�����lC�t��cc��M�ou�/u�D��sw�e�i(��*��KO�� e�d��_Dfǌ�p�$��:ܵ��O��(�:�j�i����_�l��e�Te$C���2w��xb����/��d�TϪ��]EyXF������l�6,������2��K5�8L  E<��:��K���hF6
D�Ǉ���s���TBM�SZ�<��WRFDHh
$���Zs�C�HՁk ��Ŗ���H�Y|yI�� ��3��ן�a2�udm�X�b���.���޵�O޷��+6(`�V����˨��U"��R6aDy����g�m,�;�m2c�1�y���<L���k�>S�_�ࡦ��������|�{�>��R�xK������h}cŚk+
/Z_�2)[O�w���뗭���k�h�W��j�C�H���k��HVG��@#����`�:0�7{�����H���B�V � :�K����#,Ѽ?��~� ,��%��{:F\|�%�<N�nOO��߳onݒ��W�y]�N��֧���2�����6�u�[�)�i�z,p(�Ѱ�-[9���S����v���܆OY��Y�z{��w��u�>����O�(�UW���˶��*����������;����\�4�8%y}�J� D�I�o����HD}�x�͂(Ɖ�07Fҟ��Ox��^���ɾ��쩎�VlueXe�#��!����Tl��~��71ݻ�؊X���x���)�4ģ&cʵ`��Oe�+J7�}*�1�Fc��r�r݊�XWĨ�/�Q-�ȾX� q�}}�'�{R	�yf�s?F�G�<"��b��	��ȓ���검ź�
2�	��Նz�OG ��b����Or��E� C�,�w R�*^������`��mη���'7m��wl���o����7��z�N�E�( �	/pF��B�������<�S5#�c��η9�5�s�s��O�*�'זQ�"�I��b���ɱ}�7e�Z����J+*#�|�|P)Yim�j�v���p咵O�vv�Ƹc;A}��VW\ckK�Y�������h8uBd���j��uD+����@�?��`-��:m�T�B��z
0Sw� �ݜ���S:��SNP�r�^R��41Xt`)�N�����޹c�w���e��?�X���=@��/ t����>���6@ZT���-]�h��c[�>'�U�Oմ�������ر�@�o�*�����U=17e�k�)]��,J���ʨն'w��^����r.,2�#��`&0$@7����#�;~�y�02��n8#��s��\苟��-�Dq����,��R�����љuwm|��7@��e���x�%@�+]�ڋon��݇f'�� uÚ�ֹ���[���f��S�f� ��L���V�F���S|RH�]�X[Y�@4��CN1�����pP2��Ͽ,<M=����y�"�ϔ��Y���gxBo�����d\9������Yp?�@�&p^���`�CպVͶD�>���`:�!�j?��-[~�-������֭#�5��/�g}����%��@��:�j�͎�qm���i	E��+��ˑuu.sJ�g����j0�����b�{=�(�9��^Y��{}�^��C�M>^~��v��7��ش��{v��u�[�oGV�X�u�b��;~��# S�ͧ#U�#�߽ͨ��l�D����+����'a.�Z��m�@��^ys���Ȍ��_�E�L����y}WXN?L�AXN�K�~L.�U�S��? �u��@�r:�3U6ؤ��#dr��O��exӑ7 ���7�
]�0�-[��9�~�][�|1�� T2%m=SY��S��_YF� @W�.��T9%u��^,3�1�����۹w��>���(�]IƷ�Ԥ��'F�4�O��t��K�����̈��҈\m�73��¥�� |lP�RnX��:����dU�*�8_#�ֳ{!������� �d|u\�� ��7�SN/�}�iG%�,3U)�b=��mAT��)k}:Ųշ6u=�H;h�p\GUt旴!yV�F�N<�z����2���j7�y<ID��I�<~�r3�P�}U�@D}uՖY�$𾹾n����ñUJ*̑���&��{��4>BN��)Bv�gz�}�z��ծ\�͏n��;oXie�ߤe�^U��!}U����t�����#j�@F����g�x���#gB�� Ti�y�g#T��I/@������X�e!� ¦�+Vjw՞����E����sv��7���5X�O��ïo���]+�/4m�+����V�|���ɱ0��J�+尾�� L9�ݢop�d���G�E���I��D[�~$2����)/��o6t_Tb�Z�#.���aP�<�|�~SxN?,�AXN�K��dT�#��HF�������K_8������cУ�:N?S�H~�a1���a8�3�[Q����z��X�ub�N�� ��[���Q���U��֐e[�����4z�m���qlX��|�y��^�X��?��X9m�w���,K����Y�`�E%�S{zO�w������/��xz' ��_z�5/��`l��3���������P���TM@h���Y��NO�$���t,�ߠuj�/^�ɋ=�Z6��>oK�b�b�����C;�Y���h���a�u)��*4�[	��Ha-�98�l��� U����n��^���C'L��y�J�t>%t�,�w�1'-�������~ȧ� 6��Y(ӂ5����5;��j|3�doGm�D��Sf|�g�h� ��^bS�wum���9hO��P��m�?��.~��-
��EƢ�jS।��!߱d�G����|�Q�Z�G�T#@����Z�� B��#�6�oks�	?�ӥ�_$��Ga��#:�D��;��v�sBC%�5pJ���dgK��uNZ�wϬ�,}�[���v���7�>޹{ߞ}y���ذ��m���m^��|������r]��d�-!�k�/Ӡ,_��)�c�1��:f�#3H~O�F�����@V:6r=:<�/p,遭�v�t7t�q� t�jxN?l�AXN�[JF���/d����+���U�7(a@��CTg���04�Q~�I�Q���]>���N$�����N͚��V]\���vW�+
�u�_X�������v ��]Qd,�ň�C�:/�7#f�P��	�d�:g[��dd�&#'k*k�z�y,��98����k�(��r����s.rg<2�><2]q>3�	� b䔆������n��?�<굥C�xط1�z��#ݺ-�nz����ݓ볦�Q0�\P���\3e4:)3�l�a�,/��;oڅ�޵���@"@��ln�T�pAM]o��SdP�?��S�:��U����Yy�|,d��{�L��P �}zh���̞|���[�Ʒ ƣ��9�� {W)�LSImkU��¥K��\��zv|t�m��۶�ꊽ�'lo���l����>;�R���Y��C���k���l��}��3�Ƃ��R3FBUsث�~�'F� ��A��6�'�|�vP��Gra���V=
5 ���b( &��F���C�����r5�['�WjG�s�v��v��{V[X���ڳ/n���g�荬����qme�7�=��Ϯ��R�)p�hu1F��-> � OݐVV=Y����P&�h��d�5�h�<q��]E%Ք�pŵj6��`p�>,�c���e�м?��r�����4�B�������V�ub������F���e��@��`ç8L�3#`��#;�۵��C_+F'� I]k�GG���=��/����00t�c��@��	�H X���t�2 |ػº�k�� :�y���)����/c���yd�K����s٩��t��J�w������dSRT^�:|�/�*����	S�>zx�� d��=��*��7������a��I˚; VI�P�z���W���F����]����i2��I�Z�;h��޶7�s[�q�
ͦj%Þm�o�e��?uOׇ��$P�Gy�%�0dE�Dz\�֧���s�^��eV#���Ia�S��dh��{�͗�Dnp|( B�y�2R$����~��x�];wn[G���]����֠�z��쓿�g�v墵U��ѡ��s�v�����_���_�٣'6>ط�Y�GsC~����o8��m�7
�=X��'���w�}�2��h�qO�����P�Ї�u�Θ��A�=� `lQFi*�N�����.�H�Q�o\�+���E;�ݵ��Z��s�8���$�6����ϓ�6P�پt��V��>��)�x��_ Qz�ތ�&y�~���ۋ���c�X�?��Ů�CG���S]����	�� �s:?�p��phޟ��r���f]Ԍ�R�D��~B�x0�`Gt��������{:w�����K�%@"���)JI8 H����;þ���Cv�6hu�x���x��Ӳ� ���ֺ����>����6aq� �/<VG��F�kv��㫔g'���,�$=���Y_����}o6���^�UJ�t~��ˬ�� y�gA30`Q@���!
�ȘV�����I���1q %�aT<��p p��(K7�N��1EU*i<��\���k,-��ږU��vrܶ�Y�&2dh���&uq�rź2jd�K������W�yE�]�F\Œ��v*�����v��C���O��Tߺ�����-H> Ć�,���7"�㺫��F��ҽv�� �>
�<�ݥ� ��x(C%ē�DkU>��K�>���x�`�޴���Ue;zvd�v7F�&UWm��5���#���	�lڽ/���_}m�}kZ{�fW�������?���U�c;�u�Z_'^��̺��XI�|Ҳ�g���Ha���Ɩ5�+�FU`��u0g���3B?�fE������g�q���? �?�Ț4������c�]��eϹ�ʲ����u�j���{{���_����!o!s]u]|ZQ�5��v�m�~ך��.]{C<V�L	�5��3�+w]OI\W����_8����� ��~�>�~����E_�'꣺�^�سZ�jM�?�}���u}�����{��ns��R�rzm�j����0::u���}��={��ػ�;��#�$�S�P�Ս/�`Xb���@�/�[Y\P��sJ!���
����������xg������q��a���s�*�rX#֑�\&o���ӗ{G�Y�b(w�ru[��m��%�-�(�9c��^d�O0Ѫ��J�>� "��F@����.d2��!X���S��HW�܍e�K�uY�seݧ��ͺ'jV�:�qg�7`��WH*�c:�O� H }t.���uP��7߱��S�z�=+--YO���s`-_`|��/���U���t�G�ued�,$��k�~�K\�s.\G@{�H�r^'y`-�骺8�Z�m����X��m;:;���m޸a�>x�.xS�,�΃Ƕ��I�7���p�7lc}�v�>���a�oߵ�����Xiw��U�>�6Y�l�^W�l����Q[��ª�Tϧ~+\t�*Hu�w^/�U�B��l��3�y;���NX��"p�OB(m��=yK+���S��������`T�}X�B����cz��nu�;엫[�~ݪ�]6t�ډ�>��Wu�:�����1$L��Oגz��+#����8B��e�����q��@������Ÿ�������\h^�Ы�9�0)a9���L<-��tG�����������п�6HL�X�Qtz������GVϮ�L��GFj�Dkn�잯�x�e�w5=��6v�/p�Vb�������]�� 2��7oG�19/����2<]��p4��B���|�.���U�VT�rT ��
������?T��O�(}�0nd<%�T�dU8o���G<�x��)3zL���m(>Cf��hܸp�G���E����+@��|1e(��X��arէs����l��ϥ7�۵?��]��'V?�n���Q��^�&g-{VUi>�\�@up#�	��^.2D�1N���r��!��G�������4�AR=�SK���(�>�g �������vE �-x+��َ�|y�Zw����;���,�{�=d���=�	���u����P:Q{ej�7�{�`��k+P& �h.Ȳ� ��P w$�M������DS��'�C�/q�׌w��0\����ѽ�v���UκV(�n���+6�V�\z0[jZcmݚW.9Tզ���W�s�S���0���p���܏�#s�t��~���:1|J�~E�b����Y�GG�?mll(|$�ЁYc��Ey%]>OIG9�p(a9�RG}PtN:�6#u=ǇG������Nq��
#�{���+�8�%��0��f1u����4v-T0v�x��Ny1�C��:�E&u������Q�(������X_e�Ć��v�O��?��-_�$#)C)��vʋ�C	��N���ӱ\b��4Q$i��rD>~^g����P�	%p��I�|X(98���������P�U��\��%�5b����	�V��ot�#G,  t�IdM�/}v2��>��6n�e���l�|�hMŖz��'v���?|�ߢ� �p��1��|2��V�m ��r�6�B�)�V�Fr)o��'��X�D� S�#�)~\#>�^iԭ����ꅋ`7m��_��ڧ�/nY��3+���n��W׷Y��X@��e'ag���?[�7��@VUm�$�2���;   ؁`"��C�d�%Zg����( �+uJ���!W�"Fx���&�+=�����H?��̉/Ѻ�vv��(奃���^rj\6H�q��\e����عk�l��+��Yuc]����q/��7x�v7�� #�D>Ż^jHL92��qI�"k�o���xc�7)�J���˺�����&�?|�AXN�z�k�.��:L��xvO�����6�w��0:�X���_":R��ڞ�����;\�Y�:سc^��ߐ���������S���LVB�(���%��Ii���7�t����֑A������?�� �Z7v�&��w$��K�0(�2��ag��٤�%
��2=��뀔��ۙ��ū,_T�u�SZ��Dr��'��U�b����G���=k�XK`���k������A?,��x�2ai��2}�Qh��ΠgLޖ7�l�ݷ�-]ڶbS��T��c�:��X��=ۿ}Ǟ~��=�w��3k.4���4��Z ߴ�1G@��j��I~�A�`�"�Eħ�+gi���y���a�!����wA��i���U��꺭�;oK�v�o/nݶ��o�����q�>I������G����@���ǵ l�r	|X�(cAq�pǪ=;�K�����.����߶��9]� �饬>�~D��ܧ�}dUm�V���$��ڰ;~�Gf�d��w���a��|L��:{����#p>����x]�l�_����ۚ�W����ܶɷ��c_?�0u��U�3#�p��ӟ����9re^��@U�{3KO_�#yj��������	5�ײ�=#ϩ�%?4�O�C!C�g9�p(a9�Έ����ŁBֹ��<�[�n9``|Z��O������;P��<����3:���;Lu�<�&щ�ge�iW����e��Eۑu$|��7�(�/� O��!x�QJgN_�$^���e��H��
��67m��w���̶>�)#�l��0�I��O�f�):�@9@	��,����U=�5r�:o�4������@'3F*�+뼦r�Ff��� �	0h����GO��ĳon��e��.	��v���֗m��;�6l���Xu�)�Z�֮^�쪯���t;�;�ޓ���ן��_���_X��3Y��P
�"�q�^���l@X�1iT����y;�ڗ�J(�@�3?��u�,���?%���E���.���OI��'�e�)��X����n��W�X��3�XUh�A��n��ŧw��*_���$��/~lt�H%���w�<��K?����gf+W��X:.
t���5@�W]�ˋ�����-�e	�#ǈ#<ډb���r������c=��X8�I;���P@��U�z����]{�Û�}��m;�}a������oYſ�
��{p0o��{�!��Q<�k�#�)�mfRA0�N���<�.�#��3��~
e�N�@��vlye�u�4%��l41Ӊ(ڦ������)a9�N)u<S�N��ٱ;�o�Hz^?=��Q��
��0�P*����I�Q�G�FLy��V^jZsc��V�)#�گ%�R��>k�t�ژ��#Yd����+?�0����좀GG��Dy���m�����~b��E�H4_x�Ι�Rc�{���"�b��0�n��-W�yj�/�QE:�x�������C��MɅ�!��%�����G��`J��&�
\�l�N�7���S+�Y�ݳR�n}�i�ּt�6߼f�&�=����7��ƥ��U������7maeن���l�ܽg��ܵ�/��ӯ�Z���*��������⒭ln�[��suMю�)����`Q�����ӱ	��fT�i��8�'�8�Bho�+�P ���� ��i�R`Q�>|dO��o����V8���}7�(��EpVtmj��M�On!۝]`���c���꿀�
3�[�n�a�[�����?�c[�~��kB�F:_D�V+yUn�A|蜲z����-�4�+��/��&<��s*��ǉ�B���( ƴ>�$�ֺ-]�d�7�	��go����;gv��7�s����{d��Z��d��{OG=8I׌Ҳ>pR��ڈ�Pq1�x�y��w�]���Y�	a��u��	pe�t�s�4��;Ճ�0kY�u�w�:C�K������C9��wB��D�NG���O�������O�̀B�|�(ub8(��	�:6�q�O� G@Xybo���'#b�j��mmn��Ҋ���:�3�l��)�L����P(eJ`+U�[ ���sK�V�ۑ���߶��޵�o[ck��,b|:m���@F�&�'�%A_�c"��{eH00�*=m(�%��j�+�(�����?���k�s�S�f���R%(��(#z�T��!�J	����bM�Y�[�;�����KO�+C� x�'�إ�W�&�v�t�v�>��@X��=ֶ/\�o�e�k�v�b�|�=��3{��7�{��ƻ�V:i���,;��v�?�)����To�a� Q���(�~ -rL��N�^�fQ���tS�C����4--z.xz�3n�7G<���&_n`g��bú����*l��dc������ᛛ��m�:�� p�����E�e�]�l�~����_|ㆍN|�[rx{ � �\=��]a�M�Ψ��<���/��@��E��Y�,[�p�EZ����D�(t��Wmi{۶�]�-�3�;������N�<��]ƺo���]��#3�7���}$LW��+���ˉ���e�T
��!����	@��W���q/%�9"{L1R��Q�,-���e���d9e�����Ï|)>M���á���;!:r�t���t�2�? �o��`W@�)��:(_|�uL�T�F� �D��Fc�D6J�~
p)�ڀ(����$�o=1<����v�|��펃&��bueg�P2�!�+ժ������@@c�'x�x� �;�y�U�T���Tj�lr|d���ޝ�v$]L��T~E���ӣ�]+-ӄ>���}�:���'pՋj�:��x:���A��z$ Uu`:݅�RZ�t7����
��x���C,��c��qvtj�V��=	T�S]���O����Q��=�s�}��?~fU���B��9ӊ/�=�{_}i{w�Z��1M'�Q��~,�Ǜ�a���}����%k�����$ŧ�6��E:�xtD;�nB7�*��$o��,<�!��4ڞ�,�k]�\˺�|��L�;�5�)r�P���Cme��6��ҍK�v㊝�t�ꕚ����šuOp�ذ�O9�|]�t��U�)�'ض@o��e��m�&�0 �T�Ta��4��2��Kr�1�'%�6�m%t	�D���'����/�����R������c�Tm�u^��Ӄ����}��UtO�N�p��b�N�.ܼ韵b={�Ń��RՊ�UE��y�.����z��G���CY��0��3��x����ا&���6�g�� 㞤]�ނ��;���s�ä���;!�����P����[�!��D��Q��N�Ӵ��4��GG��qYZ�� �=b��U)c�{��>a�V�G/��|O��;y<�/moغ��W���=��^mS����v�w�һo��Ң2G�6|����ۋ/>����_��7_Y������&	�W�"#=�3@������@�o*)�Kk����<��AQ@���hL0VO%�D�!/@L��O��TT��c�  kԊvR�<�+v㣛������'����_�����XY:��'�F,vU`����^Xk'�]��}���M�cc�u�qN�����r����?��n���.��ΈT��'c�8�F^Q� Q[D7�A�v���I�u6��e��^PS�lFj�M_�2��!-q��6�m��U�����u횭m����v�d/�=���O�ԲB�z��	��U;��^L�}�#[��/|��5/_���K Rd�������!y;@D�8��:���ſ����^���?���#��"ݴRxZ�Kׅ{�����T;R2�D����l��={��6�ݵF��[st:|��h���ҍk�p岃o�8�S��!�*��r+,�L&�8��>~/���Q�1:&�����雎���Nԍ*�K�p�h_m���_���M�T�����H:���9�aR�r���|GÛDl�z�>���N.:���W�����~)o��8��o�y���R`(p�м<Rg-+@���Y@{8u���{$P%��N@���+2�+vA����+�kwmO`�st��F2c[�x���ُ���w�$�0j���|����ڞ�ͯ�ŗ_�Ƀ{֒+꩹��XG`��i��
�U�E1��թcO�������Pu��۩��*�0�� }Z�ΉR)��Q��:_��YyXQa�Mz*ObԬ��Tj�lQ h�����[v��w����֨Vm��C{��7v�����1}����&Y��;;>���i]F�����	� �lm�t�8�ղ����:�̭,[��a�|M��LE9�GTb̨��
�¦�:�ŽD�S�ݏ�\�dU�7����d�C�c��ٸWm�kVb�_���7߰�~���������d��Bó������Ӷ�_�x��Y�R��J�J7���ؖ?��߸n[�>�8���{�:�s����q"��I�K��D?�$s�	����O ��UD��(8R��y�#��t��q]s���66��<O����&{{V>=�r�5Vcx���[ƫ����+>R�� F��3:����x	������n![��UP��8�C��	(��D�y�se�/Z�r��6*/�6�� �'��C&|"ߌ���0\N�����~+J]�|�@�.d�%ei��c�ad�?�/���G�&zB�Ai�|�8v9F@x��v����g�iC����;H�w��4�΃(��2hb�+l�J��:l�~���rc�n��k-6c8R�.�*#�l���+o�a+kk`�y��:�VR~J(7�v��wl��u���=��}�����e;_�_}e�ǏlA`�.�l�Ȕ��ߨ$.��5�V|�Ͼ���T����P��z@x�v�dZ��F�RF����i�0����i�)�4*�*#�r*k�0��q������, �w����<�ݳۿ���upp�k�������ic]�N���'�!}�+P�$WW�FL��X�7��t0�5��|]���m�ݷ���e�z���Y_�A���M��x�hW���#��&"mb��S7�(ң8�L�(��W]�q���8ʤ��f)�~������s���[o�9��oް�/����ןړ��k;�s�:�jGݞ�\�����ƶ䍷����Om�����XY`�M�����0J�� ��M���NO(�&��k��g�us���=_�r�*ٹ�i�+1�#���$?��ަ��K��4�b��"�b?=�[��2�RMu��X&�?�N_�F��M����v���l��%��|9_d�������'ʀ�J�?D1��tY��b�>�L��}^�ё�G�D}�W�ȏ�B�uVx�
L���W�#�$]��=�+Ź
{Y�9�!RA;�˜r��&�TP�{#L�Cܘ*��Ε�z�Ѩg��߱;��W�:��R���ud�T�i?F?�|i�ɥ�	J��"��r��N- d@���H��Sg�%)-`����Pe��v�����_Z��������5�x�]�|�.lm
|=��_}i��O}w��PO�����n��ū6h����#;�۱ӣv�?�a�XE�osX�N����Ò@�r�J6l�w����Ț�4V.�i��X	���E��:�f~�����,�FF?:u� ���c,X#���nl1dJt��":Ե��c�0���d��>�����v�+�>�=q#	��K����7��H�W|t�z#�; �d�ص49�LJ7*�i[�ku�.|�#[���Vy�.m�h�i�fͯu�+�PV�����!Cu���h�VΔ%�t�~�d �?ޔ�[���=#�HC�0ԡG���I��oK�{�����r���1b�ۮ��RK����//��{oڕ��߳�oYk�jC�������.����N����b�<?m'�$�k���� _&���O�S�l����Z�-[���G�W��D���(�rv����7iG_ߵA�c���-�qͶ~򑭾���x��}+��7}O��ZHh�s N���>�d�.g��C^��*OIr�`�=܈�h�`�7�e*��777����b�g@pH��F}�:��QF�g%�9�~S>��oE�����;��x�T���*�Q�b�g���n����4��SO���	�/M�w�M�.Q2���y���2���xx�4�,��P^����*�'X�N�Z�j�n�J�A0�/�l�����ۥk��������>yd}>��R'�86��ѯ���{|a���s�k ����a�>�����7�'��=98���UW�Wm\��h������QW�L_^7��ly�c2���G�<䑋�f�:���y	G8y�O�61���ً}�����wv�tz�`�!�BU׻�k�z5�_Y�]�&�ba�Jb������H�X��"�GRdK�ꮮ�:o]�'b[?�Ȋ��f"�N��R@KV�)E��C�����HQg��*��D"��bN�3��Ϝ*�:�ldg�p�f����7w�ѧ���gV�vm��Z�\�!��J8�׬��`��go���.|��V��M�b��ͮK�D
%,>l?��e��Q�Ԇ����Cv�eT)^?��#�uO�-�.��#���[�KO�t6���b%�zF��j?'�����w޴7�觶���VX\���{��#u�фe:�W�>��-K�!�'�]npM�qVQ��?�E8�o���c,�o<�����ۼd��W��������'�ͮ#���â��~�)a9�VDG�:����'����թ��tu��W_���s;|��Z;/|�՚��EGT�X\�'h��6�d���: ()'�<��g��'�3��) !�S<�x(��tq�.�|ˮ�|��m4���;����;�=>pUaꂵ@���ۙ:ܽ�];=��f�b�������,�a�P���=�*���媝	pM�˶�}��]�n]FD$x�6���a�YV/9p�0�O�M<(��Ia�"���A#L�dd��O�O��-�ڬ	�R��س՝򊺾�(6j�iȿ�dk�.�ƅm[Z^�?�t�6���2��b�4F��ܪ6�ܰ�l�D�~��� St������`��J�;�T�,m��$s��?§�<,�P���K���e�l@���f��%�>��6i�lt�2�J�G�?����h}�V>z������q�{���
�
���گ��笆\˙/U}�B'�W��^N'�G��_*Jig�.>++�d�
�T�yңza6_S��Ĉ�]_�z�o���w߱��m�d�=���p�-�"�_PK�r���S`T�Σ� �6��uE&�q@/���/�ך��])�xy�;��>����.������|���ʊ��	���H7O��!3�s�C����[��G�&���
�W#N�_ Ƨ��g�՟������- vt��t����e@�ϟ7�
��!�X�x���ޡE��	��(��wD�}�c�;M��4�S�i
���51"F�H�+�ť���m\+[�^��ɱ�ܽk;|^IjEj�)e`��:��}��:뚞����/Cc�G ���<�+U��w|-�
�6��5�l����'?���7l�hZ�����:q�0eG=�L��C�SڔApД�:{Z����iWM��)Mf����.6#��>�_T�]C�3�y���=;б̞k�K�\Y�ŷ�ڍ?��]z��ӃC���	���������
�U��z�m1���V>��N���55�rA�If�QY��#Mn�����QO��(��a�d<M`�1�h���!KDׅ�(�㈆�,Hb8�P<i��ʫ�S����������7;��B�f�� ��~��%���Gv����-���W�Ĺ�JV��V ̕J~J!�- �ƽ��{����퉑/��������4+/t����"w�8�c͡���@�$�:�hK[��x�-�~nuź�Hj}�g�O�qG�q�D�K�P\r^��|�py�s�9�.��2s_y[�Gr�Y�t��5�TwOC��(�{� X��t::gCצ�� ]U_+�6�}�i��N9��(;d����r��oEtt�t~�4�?��Ԕ�ꌆg-����������o}c��n��Ş=|��a-�k���d����v|�.uX0���?:���N'u<�v@Gg�t�^=�<L���y��#��P�띶�Y�����g��щ�<|⛊�<����� �ÊoJ2���!}�:�Ŋ�vc��XG���T;F�&����z&%�����v���?��₍nj͆�Ϧ^�Ä��) C�c���Q����I�#�_@���{�/�(�D�&��g�Huè0���u-7&dJ���W޼����]�b�o�a��]�a�mOnݱC�a��G���[��GWu<E�����v��?���߶��RD �����@�:H�L%�.$G�$i���P��Џ��:'o�.��_�o�?��%	�/K��2��q��"/g�#�����Nl�Y{�nշ���O>�?���޸n}]�u%el��/.0m��LI��0=�>��)��k�c&��8_ݤ��K�Eى��y�ɟ1I2$0�`IJgĊix>�c��ׇ)Բ��¢��:��C[׷#�Zd�6F�T| ��p�[�.��.��_d�� ��xוG(s��Q9��j���� �@Q���9^�2����q{��/q���)k0d}�ld�|��.rYE�����I9��":j���ި��p��>�Ƭ���W�������O��̞���6�۷�����-�X[M�����T��o�����:���K�O�G�9�J?�R���/�)��E��萋�
-VQ]�::����v��1[�����s)�_)Y�iG�R�i��+W�~nٚ��F��xFwг�:�^�lg��-�������}�z���/\���T�S2�`�T��|�O�^+��{8d�������~��ƑJ8FYRǏN��)��T6G�79Yσd�1O�+[�z�5/��K7ߵ�|���Ek�
v���}�iϿ�c�V��}���~
֓�Z*�'�,�s����� ���{V �(�	|UKl}���F3�Y�p�~X�h��+,�kM�j�?����ֵ!?1��.cṔfʛ��s�\�=��)�ϴ��r���X|~ɯ�ə�C[~�M���e��7�[�Q0F��C��Z�wُ�JA�\�L�h���k�`?���6D\ �HOۈk�uDv�Y�΃����LK�<)�e��e1,	=B�LeC�;SY�~C��_X�U��������b˵f�?E��<"���z�'�)��:S�\ڹ�u%E��?���>�PFD�42��q>�߀8*���C�����q���D� G�n�a9�~S�vdN��l��Z.F z,�n�V8>������h����m�eK��u��.wh��:H�`ԁ�7�l���l�G���ZsC����:u0C�3�u�Լ�z��	��E����4�f�4��Ț�HGv$�y�F4O鬻a]U��~�=��/�������Ͽ4�a�ᾯ�Oj��|ʒ��7�mku����N���N_����
�"rЁ�Qy���e��������}���VWlܨ�(\Q��:��Bnn.3��^�W� �3����#13"���e\ߌ<�\��p�ʣ�e]��T24�t,#���QadF��Om(����S;��۹}�*�U��M���e�O���k�ָ�mo~��F���r3�*c�
��Q�lb�F��%3�j�"M� R7������qԉZ���)��Wf�U�Х�NR��K��~�2P�N��f	]����L��&�pW���yC��t��]k��Y����{���E�1r*䆖��� f��0�zR�x�p훇�C$]q|J/$7~x%`q��:�"�y����*�יS�u����� �)����Jo;�w�6:�1"躤\9����5pYyrh� Z���:^d�H;�)��˙��< @�TӞ�a�یγ�*d�v��QX8Ԯv�v�ߔE�ҳ�<�u���R��j������Gg���/��K�\�$�|�ۘ��\~��/��~)a9�vԧ3P'T�X��(����;�������O��k��<ꣁ�Q�GZބ��v�"���m������G����VY^7v�f�pf����G��13"<��E�g"������#����E:>�C�M%�����=��_���ۻ{�7"�*�Ԩ�"�Z��&�w��ۭ���<{b��S�Y�o��̮�u0F��]��{���=[|C��d�y�����M?˒��g�S�:_��b��C��B_nв���8�cbṜw�%C�ytQ��W�=S�z��<;�c>K$�u��_Y����.�U(�T�֖��dH�.��;��ʵ+vQ���m�ܦ���鱦F:���,���~%�UaJXG>��J7�:e�΅F����S/���$N�ݐ �&R9���!t��g���* �QR�"sǝ��$��ډO�ZӉX2*(\fDU��*�M^ل��Vtu�}��7=Qv" ��.�����'Jm�?�)�W菺�;�;�J�u�$Ӱ d!1�!�{�(�A��"W���\+����(���9o9Σ0$�f{���]��N �Q�o�����м^`��7�$�C	琏�I�{9�I���-K�A��M9)�[�~��,�#��G�"!,�g�>������-�+N�O�^%�q���XN���OG��[R�|C�
EAX������꿱���_�u����\��<Fr��F������y�NJFgR�YU@���B�d�K��:<��D).:�Y��ߏ��7Q�����X�tʹOG৓剕�3F��:��₯c;�m"���s���u���M���[vq��u������v�=��Y�r�^ߧp��G��] [۴|ho����[oY_�:���'��(�j"+�ƥY�9yT�'��?a��pм~���̹x
��y�t$*o����8�q᭿�GO���=;y���G6����VYα���ҏ�@�vn�z 1Fg���+�/
P&�a�y�
G@��Q;���1�����4I��M)�'	.�{#��Wd �Ў�K$�A�)d����	C�3�Qg�l��!�]a�!�Sz��#�:�9;�\\F��N۵G����%��\qd�2~Q�����Q/�(6��[I\&��	i<}VX*"mK��Y��#�8 >�<og8i���5����6�3��QΧ?�s��(�$�\�w=��.�x� � ��+0�H�>��9�a '�WG8 ��J>�ͧ��r�:��Y��������s������[�R���V�������'������������# Xy��C���e�0:�<?�Sp�۷R�a���W��Mu&a|�h :�0�q>����:!:��aA)�Ȭ�L`�����,���aᕏ��>Ƣް��UVVl��U���;v��wl��y������v�/m{��������T�˃��u��f��Kv�O���n�o�i�zMq��$���c�K���XQ/����iR�L�-Q��7S�)�r��f�{����$KE�4����7;�WҎ1"26�lQcd�O@=}f��߶�٩pv�:Ñt)��V._�s`����/m��I������M�,Ԗ���2j�Q5�+�ŨF̍������ ��!s�H3�H���69�S��Y��8s<��E7Y����,�@e1B��`���S�E	�	���;++]'��#r9�Wu�(K2%��Q���Oc���G�<��D��s�"�(�	���T`�p�(:�G���qd��m@������#����H�|�y=]���Ku^V��'�7~:"O��<\�{-����8��>��h��K ����^YSɾw|�>ēr>�;q��D)|>>��?�ӑ9�Vԕ㉽|ֲz�k���_����G��NnM�d��S��O�-����Xg2�o �o.إ>���?��wޖ1�d��%+2��?_C��T:�i�D�o"���S3O������ߧ"H�d��*������c�6�����XMu)	lF}{����\뫯���ܲѡ _`�xFU���}���m���֟���ϝ�OYp]`:JV'�	7�22�Q,+�[fbR��lNi���Q�0�E#�	'�4��7`AI����m�l�v0�
�W�<*{Y��������Ϳ���s������Y\۰����?������ٹMԛ6��"aQ>��n���56���"�f���<��1BV��� 2`�hj;ӑ��[�����З�i����F��i@�/��S�Q�LO��U�듖�v���:1�]��}�C	���=:p#�H��_T���偀�
k�h��D���$98Ɣ'�:�#u��$g����s
�����?'�I��4�G�|*T��?�֣����A֡�7�Q���r���A���4Ņi`���ewP.0F�=���\��0x��D��!����z��)�4�L�AX`ԍ,�N�/�l�����:#M�w�3B�|�v��_�E��U
>1Z��w����K�HXNNѵ�������ޑ����������:=���O����K[Sg���d�n��D}�/����6��(W��>�%WY߲7߷?��]������u���%:�Dt6t0�Ir�2J�O2.����#���4	���f;�x����m%X�_ �Z��?�7����_���;V�|t�[����g
++V�\�y��?��.��'�z�-�>�&�$9�'��1A���^��u�� �|�iI�t���Co��y^��0ȍ)y>=��H@�$����ȖF<�0�p�8�lԭ��`�j��Ol��7[]���߲k?��]��#+omZ�Q�j�I&/׷���R�߷t`�
f� S���Dz��"�K�Q�-��|�.����DQ/��~����1k30%e�������1x��	U��WJ���/)��/�(P�qb�]7����Q|v��D���v�UI��C�K����?g� ��kg���8�=w�C���b��q��A�v�%P����O=9"q���,U���1�������e�J����⣲^V ����.s\w�i����F�J �tA��T'���"�!����b�����V��i���E��w��L��~(	��	#���:��3a�8�)ֻF���:����l�����9���KV���wh�G���}Y�:0�Wm�;�Tl��d["��S[�qՊk�6`W�:��+}��F����D�b}!��� �z:G�?ي8��2u^�׍����75�"#:K��9�T�ޮ+�/����Z�G�m�?��O��ޣ�Vj�hϤOY�z�ա6��	���l��wl����8�!��P]f���O9�!�S:ן�,�����BN7"�22#"�Dra]~���|�0��di�T�"  ��^�(�|��˓F ������}}�5�W��;oۍ���*�t�*�'��e���?�9���y%(*R���g�7x�B� ڱ��_
�8���ۜ_#2���+(�S�����'�����,Qg�e��t�U��yD&B�����˛r��|����*عy4�c�#de�N D����q'�E&#O`�U�A�j��r��<L��GM�)�>#���s�#��",ڗ�F���/B�{>�{Vmϗ��\vgM�y ��F�~�Ei�Sg0��8�_�%���Zr�k+9�s�+r1�Ś0 �.v��	�s(�&VWW�ƍ���@��"�7m2Յ#rrLa!w�aN�w�AXNN��ݽ
�h�4x��:�	�J������G�[������s6���َ��Zw�ؿ	�IE�t_��~�g��5�~�}������oڰY���|4C��O9�D�c���T�:"?r��w8�EG����^%:( <Rg�&���a!�OF$�T�S_(k�tl�t����v�/��5���vr�,�.�@n�д�kWm�������+V^]�r`�(A��j��vQ��%b4 ]L���d��E�t�/F��/#!�H�c��Ξ=Q���8�IS*쓦��F���9}4��(/�.�&��ٵ'ϟ[E:پr�ʍ:�2�|T|b��gQۓ]���u	I��'�M���y�n_	`�j7�t����๺�@Q����r��J�<�
�z��E
S w�&K�||�2R�s�A��~��9�O�Iq�aP�M��1(�k�X��2���Hb(��S�\lـ�G��I��T��/�0
�ߣ� ��?��`�}</@��޸W^�_�q_o�	<%^3
��lS�O���+z���S��ĥ2�0d���%[]��s��d�j���WΟ?oo����E=8F= ��K������������DG���֦���1�7?��:�G_|n����c�R��J�k�����'�srf�ӎ���g�Y�1*N�L�k�а�҂���]g��7���b��5����zz��̐�&
��	2:��|R8Dg�j�ĹwVj��J���d�����Q�`#R�,	^VHi����`|�����ɽ�v��e���k�<{�o��T~}k��n\�s�g>�i͋��3M=���aLCq���\ɔꒈp����eV�w�d'}��c�t�������e'݄,�at0*�9���[6rIk��2Ň�qCnX+(��� ݱ��ժx�U&k�8Wپ�ߍcF.7�!��Ȍ\��)o�y�Mz��:��z���8��2�4i$5M�ɗ��?��P2�Q&��˚] g�ťp/���q-����7:��&��� E�yD�o�C�w�DpFY�_Bf����]�Ε�Y!/q$���o���J�q�<���KG�?n�`��$9�����5Hz�2�~���?��Y� TJI��o�$���(Q�>xEڗ��y>��~(.bO/�&i��7x��{.ʃ����L�Ok�R��/d���w#��>oׯ_s=�����8�_��o�_�R�r�~R�&,�)�1p�Fיݸ:�G�쀪�O��/����6�_��7�ݽc���6�Sd�}_��z\�����Y\��:�Kd�~�[�m�//X�$�B'�ը�)ӱ+�53|��7��э���0�ƧΈ�W])�[� ��c��QL@$QF��U����U��������p`��-����m���za�:|kQ&�X�ZE ��`����9erz�Y'�DN	C�ei^�,/��'�%���Q�����:w(�G(d�O���\F?a�FT��:)l �6�Vl"���0xXr�W�y��;/Z��r$�zqT��!�G��6;��r�2�,<KC}���T6.8�U_��/�c��tv}  Dŵ� Q&/yi�΃c���)�3��R�~>�Fz\����Wʛ�t�d�� `ԓ����*�����>g��x�����\V�'\ &J��=m���K��E��t�	T�0rN�"�d�<��(O�3�Y�8��<����y�
��6&��? ���:F9�G�|�O�ʧ6Cx�T1�V����2��v|�^>��J�!�wQ*3����J9�iJ�غe���nZ�)t�1����s��_�kk=yl��#{��Wvp<}n�����7��<�vW*6��mm�*oܰs?�Į~�
��ukß�WO~�#�f�w�"u�^�����A ���N�4Z�N?�A�y����+뤒����s>�c:��yVy��y�D}u>��I�m�Ŧm��������[oZc��ud�NՉJ�%��b}�Ai��DM��Ma����Y|�`䆟�Q��|�k�K��_�ů�˝��s%�.�%y}$B ��?>Gs�� ��c2�3��p>
���+2����n��Ϯm�3⾛���hN�0婣�@y8�)�"�̗�KE���d�3�K
�e������r�1ˎӬ���U
����W���{V�\�� V����#-2RJ\{��=�4Y�$v�'��L.�pT����'F������O�y[��z�0���"�I2�K�hCѧ��'<�י��k&S|�E^(}�+��i���AQF�e%���q<�D��Ǵ�Pq|q���C��~�4�����tF��C��r=�������Ȝ�����D��͢`>	�{����ё}�We��ܶ��S{��_���s�=~f�^�:L5�6Pg2��|������^=o�g[7߷s/�H��Hu���<UN���h�f��藞 y�|�ՃL;�tL ,u:�8�8~sQj��͓;�ީe|q������y��F�y��و�����>U�w�o��v�䉝u����fo\����1�$�TR�{b��P��O����������7�.%=�L�s��#�u'���'|��p>�>�N<h�9;=�?fA#,x(�Ee"=�k���H���Հ�a�^v@��^X\W��#��#?4S����H��,	e:��9	J�1��2�j�� ���P�dF��%�2��s����S' $W�ڟ�� Tj��k�>�"p��Fg�5���\N�+N>O��!d�"���:QwO`�(�GJٚ%��X�)�ܛ�9J�+�DȘ�A�%��ٽ�f#��3C��<F�����+}S����g<",��<���rYE�!A$�|��7�,��ʏ�T��x��Q�>�)}#w�޴7�|����l{!�:{����C�S}8On><��� ,''uw�1���ρ$ ��f	O����>���;6`o����?�g־����@��U�����juk^ܶ�o�ƻ׬r���6��Z�{�h�w���bg:sv��[�t��]D����������(�;a�%:�,.��O��T����3��%:��&Ż5�E����ST�֡��PmH���1��f������P~�m2��cF�MGD�ċ2�O�Q�K7�,^�(����q�:sA���ם�EB���23��s�����O��z)��Z�(1dG(tP�:�G
Һ_�C�y��k���t�����BWjo��>���d��?�Q?䖌D��-V�;�)���l��nLE�}]/���VvF�w=$v9E��� ��_a,�O���r~�kJ��y�B⅑���h�q�t \�b=���`%ЉmM���G��E\Oډ_O�R�#�
�*��=�t�hL�Q�),(�����E=#�DE�*)���9��Ґ�ӌ���}�~�H��1��)/�����5	>���zݾ ؚ��۾�+�,^������.�IG�Kr{�A),��=�ZFN?x�n��|{:����}��y�L�z"�V�Q�;�9<:�(�@1l��QXys��}�]��O�ʟ���|𞕷7�_.���㽬��_YO��y%O�t�� 5�p�7!yRT�3߹�N$M	9)�}�iJ��s!D��Q2�q���'S�.[�g�G1����G��_K��f�li�&���H�G+}�Q_+�f&ԁ��>A���Q��H�9ӝ��ͳ�:V(x�ѳn$䦺L}z��ғ�4F�8�ťx?�wq�Ӈg�p�uv]���E�q��g��*�)�;t�,��B6Wf&����)ɛ'R�Lw�����xey���C��|�>Y�0�P:ǫ4�h�:��M[�������(���3y�{�k�C����du���>
�4��}� ����%`����Z��׀�"_C��CV1�FE�-���cN��8%O�M�uI�)k[P♀<�����t>O��8q>�O���zN��H�8�zv�L�3�Xg�2�7�%d��a�F��_�A���8<:�'O+���d �]��9��T��u���^��br��I:0�qs��[�������-..xg�ƛ,D]^Y��:��:����U����l��S���Gּx�z�~���I�F��Nw�_NG �C��uN'�!.gt8�SI���)��%�t1�=����ꜧC�</x���O���G27���RN��;iՑNTi�:�4�`rz�'\9g�æ�G���AG���
�&'�Cܠ&6~�w ���� �D�N���Q��˚�OJ:Ђ!�;�����	<S^L�0�z	>��P�"u�X9t���|�lr���S��A�&=�M������n�>�ق'�8���SN�&����r����@y��#�jģ�Vb4Heш�W<��lŹ*�t�~�w�L�G\ȍ��ZD�Y�o��N�����~�ݑ֯1@ArV$gE1�/鼨��x����؞�ݐ��ċ+������%��H��G�uOL&'��=�K�:�FD��y�A8Rq>O��3�hGqͣ-�7b'��R��~҄\��SQ=rvO��TV�Y������z��-4��M{�bǞ<y��0z��y\re�t͡�w������l9�$���@ō�@<���u�28z:cde�ƁJS�T���h-u����U�^���S{�����{��U66�_([,4葁�O��ձmŠ4�~Q�MǑ¼R��Q	��HF�4��,�$p��I�*�S�+�Ҩ���F����+���A9ZB������^+V�6 �-K���m�N�/0�ki�G ��6
r?��H�QGu�J ������(�.;q��B�
��-��~:�K'��Rx����c��[�:���1i�jG��#l��\��E���Vq��wJ$?uvPN L�ȷnPP �YHF7c5�.��G]��D"��`���B�1�K���O�J��VX8"���E��O����F�����B�{�͈��z%~/��ʜ�q���e�TX�c�a�J]��@m��6ݷj�`U�+qJ��t��!���rT���"�ۡ	Ja!ez�t�Nn��%z�<��a��<�<s�M ��{�<��vM:b�Om1M���8���HexfQ�w>ܣ�\:�������m,�-o������A�j���pמ<{�0�H�c��|Qj��-�w�������=JN9�#�Mϑ���[�n���>��`ȢRf$�]�C�[[V]_��k��ҏ?�K?��j�m�T\��NM��T���o�!vu"|xתE���c��}Qk�A�\u�PY<9{�`:|:i��:�y�/�P��Hgq6z�ͧ��N*��S���OCp�h9�K? F V�jd��c�^|��I]���r���4�n:��x��12�qOF�:�N5��V���^���r&r�$�(��y�3�1R8��_�9(o��������G�
��FK5�C��|G��Ob������>�>�7?�y=NjF���Jq8t�S��
]G�!�����TF/�G�Ѝ�4�4� xCɀ�5��8�)�D�z��c￟$;�<OP��{p�� 	���]�ffwENN���ٽ_F����ݝ�E�g	 yfp�,"����Sw���g�zj�*���QSSUc��ٳ'7�D���u��&�:�w�_�&P8��L�����9����~�m>����8�� ���a&ë%���̗��t׈fѧ��m��0�\��G��D�W�d"m2\��Я4���$���&ʓN�^�O�)h <��O]��*j����h�P^C���V�YE���u�H�|����bcG;��O�����O� � ـ7��'�'q��/�o����:��i���Z���_Ƈ}-FX���`�7�ԉ϶���ƽ�_y»|�F\}�ո�����_�7�мf���r�c�t�A�YA~�C�b Ql�O�I��v%6�qard��_�'m��q��̀����� y��%y�N�����_�GF$+X��p�%�q����l3��#���M^�A&���a��Iߧ�J�k}Y.@����(c�	�	,)Gx�#2)s�n�>
���!�x���ʳ��I�8�N���fy�,��:}��X�80�۰���8Ё.񦟆�_��oc�|��>��
�ɇ�^�S�ӑ i͊ێh[NӖS%����V��.b��jM�7dMG�9̲��/���L2��T���-�2���߳����Y�)iփ�02�/��9�?+J�<�_&�6놝+��~����������{�8w��bf��/���ZL�-���rL���qk�G��D��.�*�h_��K���*,����C_��bh$4O��xh�^� ���퀮���Pix-�u��E�:�6���QZS��'Y�-�F�4�W���/��r4���m�ig&g<�8*飹��M� yN�Y��z�� �$=�P��m�˽^/�W��W�#YY9C�"\d��Y�丑C��}�wH87����u�	��î?"|������<���͹�j��?؋͇�c� �䕫����Ї�����>ЀA��;qт���*�9Yj�ȑf4 ����i�@���,��y��G���a��`� ��x᧸*���;�^��ifI�d�_C�4HUҨ���=���^Sz3��imd`��%���f0�͕'e����YM�g<ԟ�%�#�8�U~לH��1��8JN�2YY��	('����4qFIލ(G���#Sv����fWX�,�k���0�o��,�`��C�ZX-VP���|����MМU<͉�]�Eg3g��&��F@ry�6O S훬����!(�\#8=�%5>���S9��_���g6j^�mW�|B�ڊ6��gY���ta�͋'Cw���t ׋�/����e�y'Z�������t,\��^���_��W^����苯��,����"���I����YE��A��*}�Ϧn�+�
�!>�з�h��Fy�9}�Uz�?�4���1Q ��	��P�t��e"^��B��<���x�q`j��O����,� ^��1G��g�T�Q��(�p�#o@(#/]�/�.�ؔ������������J�C�ƙ�9��7���'
��t�ꠏ=��>���������{j"�9����/��Wc�Ӝ=HhR:w~�,T�˩	a<��5���R�'�bo�&�|1�2��ǃj����7�Lȸ����@�'���ʛ�6�\p��2r�-�Ɉt��KfLԔ��1|��r�arg@�����fC*��������v�Sͺ�}L��C3�hM�*�����/I[q�	�5�����K��
0甁l ]4FA9��W�y�,��v�Jw�4�E&͌��2R�ʮk��a�
F��T~��$�p�gmib�9���.�z�K��-O���/|�rs`��<%GUvB�HV~������!���w��%*Kg�R�f�����?&bDT�Z�Aê�4pNc�ޝ����>y�͍�����`?��;��݋�ޡ�����=߱1�.f����o_<�WAK�6LY|w�u*2� yF�G`y��|Z�3�otc�&��� �cE�0�&QP��2�9�8t�tA�9�#����w�3/u M�;���;N@ �����M��$o	g�����:��k{�F��@�*"�&cw87��������xy=��p?��c��8��4�Ί��@΃8����<�qg�@�ż�<q�,�g������ЯxCF�i���>�a̫\��cqN���,8?� ����ysV��Z�(1����
	99�'/� �8����ӟyi����$�k�(H��)�nưarg�+I��dL��#���H�&2R��X���\��Fa ��6��f������'�E5q��Q�h���*_�G�!g$7�Ϩ�\�*��^%�&y��iV����K�E��K��߳@�5>�o@ e��@�&|��ZFB�7�8�m,填9~�f�˛HK?
@�T��ê��OK���``� L@���Ҟ���v�Dws3f���!{o�r'
w����v��8�iy��,ކ��H��w�E�|1�HT��s�0y]��j'���%k�'Tު?�rlS��3��)��!$Yahh�yH�cCO�B�	ޜf9�1F���5���'��)w����Ӓ���Y6�a �$��ͭXZZ���|Jf]7@E�Z��q�����s#�O��逻�;�����Ύ�¡��/�G��K�B�����]H��� �F��� �&�'pe��3Id���U��(I��'��pGd�_�Ϸ �����9.�}�.��4�(P�o����&��4�n�x�#씄�{�81��Oٓ0*��7��BvOQS8�g����3�>�-�B~�,688��	�!-W����1O���i�����;�|��q�S/E٠i�ND�yr�q(�v����]Pi��I �1���F�x�KP�&'���HFY|�K	q&��DM��[�2Z�<����#?��T�$#�Ic��G� >��g<.����O*>���
W���Qi��β/H�C�� ��+}�rN���c'�@���J~�Xh���t?4��?و������pm�jp����������h��]Y�*B��I�'�1��T�"]m�ܔ_�m&��Mx?��D�A@�6�LO��R���D���t�����8���~ĤK�4��i�!G�'�7�(ܤ��Iȸ�c^cS�,�k�ztt++�1??o]��r�����P2��΍�?Q�� ���0>�������Fw��`Lxt�2>�6X�< ��@�9�|�3x��_р&>&�I~�ipz��!��Rt�ݢ]�\�>Wd��L��t.��r� 9*G�L�'g�'<N+��dm&�M���IYLϱ�7׆�e�Wĸ���q�rp�?�,�p��!J� �Y���v�����٥A7é��Ks�\�h� �OC����Y9�x�~(��$���/�NH��:VA�AF�s�U�0d���Ĵг~7�t��y_�]����N�U��1ɉ�B������ QB�*��&�����?�X�#�iAL�+�ڱe�,]�}���7؈���+e+��32�ZÁdՍ�{��X?^[7`~�*��i�d����M�Ӻ)k/-Ew؏#�S2`��EGv���z�.]�9�	���h��*�����%یEl�+�`�=��Oť.$��j+�0p�j��'�2�����������VꞫ�Zb�*_>�Ͷ��)P�y�n�&�'�UNB�e=��e7^�ȶ˞5�	�A���^���U�[�E����z,�*���s��	�F�5d�ˁ����9�`������?�ͭ�h�gu��ې�/'W���2~3�;���46��	+�������rd��A�	dj��PFY~S���N��jb�����E�t�<�+�ף�����(�GS��k��@�r�7 �G��
$?Ѐ?V]�� ^�X���ϑ�3�c 8Д/�XN�N�:N<����������J�玤o�*�;�1��u>�����IㄸL+:�L9��������/�.�t�5\u_@$3���� y�/�d\��������F�l���V�>�ޣ'qrp�s�hae���dI�;�1�IZ���W�¾;;�p�b�$o#�K���o���Q��w�&��V��I���H'
�"V�6Ӛ�A>��n7Ny���X�w�?մZ�b_76�s��z)�/^�ٕ��^_���Wbؚэ�A���)g�I�yasW�Ǽ���)_ƀ2�����a�a� �7�NB�/X?���6J�Sa�<A��Li�n�n��~��9�4������6�e}�9����������J�˒њ�1"t���DزߟFc� �၌c�-/���#c"x<��������s���s#����ߝ��~D����'�'�>�A3'E&-�t|�Lq�ֵ5�9[�_c4(?���թ�7���<�x܁��gpˍӤ�@�>�_?�����3��tr`��ũ��C�a��܉���$>e9�+�&� ��yIS�	��gUХ�g0�����7e
�*���O͎.���pJ���fNMz�v�m9|������:@gTN�O��)=dp���v)����l�[�&(\˩��	�v��\�h�7���l�8c4t��h��z0�1�6������~�_~�;��޻������o��3��؉�Ź\���u�<��}"MՉF"��҂��(�3m���I 煮	 �tL7[t�ө��2�f��::��ى{��6���8�މ�Օh��Ǵ�1&u�0�w��<���ƫ�Ƣ�������ߏ��JG�a�v!�����*]�u#&&`c>G}Х<-_Ƀ���a2<³�,>Y��º8M >z�?�7d���ζ�0*�!N�a�KI���Se�?7�X��@^h��cq�Kn��G��4��� �m���\���y;��e&n��Ե��ŝÿ�a��C�ʠ;)�����~�����CX=A	�4���+�;0a9h���<�4���	*f��%;��&ੀ�0|�\�����r�����l�y�_\��<�LG�܇5i �^
���O��1H6q5��D;�KH�D��0&B�2������CR3A�o���.�0閣��y�6�hr��T��G7��=��h(���k�*f��;�T��� @�ɳCΓx6���-f�Ra��CR.���k�6�d�SN(��Gv�(S�X��<�IU� S*�B>�4��ů���W1�h3�ᓘ�܎ݻwc���������b��x��aቒ�u���L�'�"��^�A#C�
I!}r�O���ڠEg����>'e�CS�vA)w�?�����������)v�܍������ta]�Ӣ�E[7Q������C�5j����e�,t�{|�;�<�9��5�W�c���h/��@�v�Ý��]�*!�����O�k��%�ӀƲ��27:�Q�xU�7t���<���/��7��ɲ�,��5a4�������ʟ�~x��d��1�4��7â�0Ŕʈsߒ����=�+��>瑰�Vz��1_	��ˆ�J�~�pn��Q�N�@��߽{��w�q��q�㩣7C	����=(Te�ˁ����?����P<�q83���&�K�;�mxβs �@�
'Mx���s���=9�=WW�ř^�\��Q�Ⲭ�<��^�o�s�] >�2��ryD@�p&����t���M8�B�t?���kG�&O6gs�����{wf���W���
��D��W��k�ɪ���G&|	U�q?��Um�,kl��?���f0F�2a���r�G���Q=x��1'��tO:�	;���(�XAR1��v,�/H]�`�"��w�r�R�$Ϗ�3汑�����D��ՠNB��h�ˣ~A]뚓,u�h�W�0N�Gq$���/~��~+Jo�Ɓ�̹ՕX\_��ď[�����ya��l�2��DgY���6���q��@���V�-�ƒ��kq"\���']%�W����6!s�3m2���˶�8�S�Q��C�s>�k�(q�o�ț��
F��\�S�����x��.���q�0�>C\q�f�0�<��.#��q胷��7ܽ?luպ`:"/�m�}��8��o�F�1�#��Hթp[�[6�؀��.���$µR����·����~��E�CÃ��Y':v(��d�/(>XUxz#K�b�3�Njh��e$᜷q6ڜ!a��=�5�H��Ɛm�a孉��1����ܨ$5�0��{�5�b�Z��2�1�����<�4C=�^�2.f��������`?fEo��BԵ������JB���� ~c܄��y��xSS2zfRH=f�1�����4�#o>b�Ɋ�Q��N��������.Hr���� b�ⷶ��wR�cqF��Od|{�8�܎͝�8�Qu��X�!&�~���[���.8��-<����ǵ�j��#=�#M� Rw���z4��?uJ(q�f�ů�ǳ��x���b�Ϣ�d+�=�鎓�ca./]���e���p?6��e|��_ơ����������W_G��n�����i϶;������q����]Z�A��}g=��ӕ7%��|*����hdl����1@�aR_�0M9�$1��(Oq�W���V��,���J���:o�@��������h����c=8.��6����Q$����P$���*h�|�P��r,-/Y^pl�)c�;�m�9�����#��'��#����ۏ������luP���y`B�#cP���@�AP��y�`̻����6����W06T�@���'S2��*�4,r�H��lf��ie4a�$�G!A�6 �̺�w>�ᡡGZ�����AY	�� �8L����}u�7��S�$��
�8ЄX�N��%�0
Xى�=�\�}}'6?�"�Y�?x��GOl�2Ffb�=�)6�B{�d����ю���8 �̓�\��A��ʤhC��4�1kh�fR��&٨&�q9�ٜ�N��(������.���0+K%Ǡ݊V�-�C�e��P9��	>L�鴣/㌷$�h�D�י��~�BL��N�P�g9�fe���b(�/�lO;�����#θ�[��)|�Հ}�'}�G�X����< <o<�#������}�-Ɇ5hMGG��s7b���8���廿���?c���1|�$�>���n��{��}�w���1�����Wb���h_X��?��n߉�΂Ϯ:�U}ӝ0nř�DF�8D��C
�|7*^1��+���������IPO�f�c�=o��]�ur�焒V�Qee�� �$/��1vҮ�r��4h�_���r\��k�&��E��5�����*|4
"S��8�ߗ��f�h������q����s#� ��& ;��xD��I���������xW7�s����Pw��̄������Թ�
�8����/�y�EZ|�.�L:���*OA>nʼ�˩��THő#Ͽ�@�҄�1��!{[�q���m��Ǒ��M��q�a>�k
����� [)U��H([9U�rjxR�(�C��'�?��a~f���M̍�j �jo�#ι��K�,Ti����fZ��?�;2�{����x������wc�ӏb�4!�{����8=8��&T���Ι�ag�-��8�o�bб
�<Z�0N���$�kB�Ա�RW˪�L#��H��0:ǯ����]_8�k�;�?�W�� ��k����8�ٌ���҄(w�Il(�s^my�Պݐ�Hƽ�����EY�� Fw� g[q|��BN�X�_�Y���9�8�����`H�_�rȝ0�ܠ 1�ŏ����i�I!�O����/h�U�jc|����F�x?�dLmݻ��2*Ϣ�*��z\z�ո|��h/��qo���x�l��f�Շbw?N����Cs�cp���������Ջ��vA�Y�ݾ_��/b��(^��\,�/EOF��bv�Ӳ�NгXC��a��a�4BsͶ�� ��Q���-��FKC����Z)ö�%��梚~�?��,��̧ ����S]S��!�?��?�C.�5c������7�Ѕ��Vfop%�p�G1"��'d~�?F�ȉ�Γg��'~��h#~�������#���R�����4���_�򗱹��;��'�~���d�?5D�V��ܫ�����'�A��Tj`�2��zi�*2�A4Lʠ�q鱁�7���h~` N�CC�h��اs�D�=r���gp4�2��L����4W�yuCt�����C(��f�\���7G_(&ț�f9����0Ip>������dG{1��D1�6(
KN��	�o=ڌݯ�ģ�ߏ��>���n,���V��Qvbwk;v�v�7hjq!�d��Oo�}�5y�/&�HO'�R�����a��&�6SiD���?��Gcd���8�����W٧-�Ե#�,��
�W��66�߉���X[[�2>�}��N����� �]]��_#n��Z\����m�H���ȳ�d�N��bz~A��1�$z�$QOܮ�v�:�
S�:"N��
��8�(��/9hCφ�&W2Ջ$�נ3j,Х��gZ������G���S����B\|�Ÿ��w��[�'�h����;ױ��jg����nں"�J��1:����qí�>ي�����؋��B,]� Txm)�9V��!��X��%����E�H�7� 0��Q�X����*O��Mr>�N�-�	']g6C��QJp�GM�B2P<�栉'�|~*H�υ�yLh�c8� ����9���E}0�c��T^��z|t�6�J{�x��Kŧ�ȸ/�̎���8q=��?�a�@�qǕ{_�ݻw��nG��v�oA5xyW�`�}�h������tH f�I��/�(��������5��{S������A��t8 o�Mb�xS��S���=��0��uZ��坖�|���a�pd'�\!��HJ�������<Y�x�f�O�T\Ə�l0��A%��F�_�π�	�v6Є
�^����3�O ��LKF���ɇ�g4�k�D��W�݃X���A�~ߺ����f;q���ԧ���L��]�b̒M �M����=~r��d���F�4��9)d��٦Hκ*}@���O�g���8'~�O6����W�S�c������/A�{2��pu_~�e�o�L輌�vG���P��^Ʃ��i]���j��^�օ��ǁڗV��{��He��;m_8�[7�2�R��i���䠅��'Y�ndO�+[�X[
�`�J��=َރ�8}�%���Y-�t!Vn݌�׼?���؜~�0��xr�n�rt�he�� w	�-����a�d�"RW�;Ĉ�ߏ���,��%��a�i��X������B�W�bld�����9Sʰ(�4顓�2\��KBy�g�5�Ζ��D����>����x�I>�*�,�/��kB�ϱ7y�X�o]�d�4�t��e|��?�7�������\���1|��%��4 }��
<�s�87��hA�E��o�E|��G6����< Ѓ�Tt+:�'�f���[�>��2�㛰�_�un`�kv�I�&Ϸ�{�n�ȁΣ� '!�+XLr2�8��$���&cM�k��\��J��\�Ct�ͺ��*y)�V�<��<~L@��*���r��0��4�\"�P�{"�[u#R�W���ᱠ'EYIɟ��q
�4+24�!.Ȩ������8�܎��}r�Lw�G�Q؏i9��!�Rg.:2H��<���#8'i�^@� m���'�4��WE ��X�ƐC^_	��IuT�5����V̫�f��c������G����>��I�|z��0���֔t4��6���O��[�0�t�]�|!�$dw'�p98�VO{�.\���c��%?������LcK�х��oR?U�����Z	�Kփ��_=�7�	�1lG&�[���������ц��S�+��ܵ�_]ʕ_�����/o�΃ѕ�Sj<~�E>�Ow�
q����f�=w�#�zJHw���rV���-zI+'�1�L�S�w��8��/4Bb�����O�+V�џ�T��w�?�qY6iy�z�<���m��e��K����d�R\�ep�7�Y�U�/��MQ�ǥ!�aƣLK��1=D����uc}m}t�Pr�/�������s�o�s#�����Ǐǯ�k�����`lh0!��D.���w���'�7@]�����$oz2�����&��끠���hh�Z�c]��� �Tt�fd�-@O�ͩ&ݖ�<>���d��n\�'�^�|����Ƽre���<�1 �ct��=����2�̩���e�4�s�6r-���ٸ&R&�"Y�p`��a�B�;��}:�p�=C�[����������y�S�!�2�P9�Ě�,!M��SGr����uK�H{uE�Z�[�2y2`���CM~b�2�2�5'C��zJ��������7y�]qi��^Kw�!�8\#������dc#n����#����a!�kzA�{��oK�ì&�Ç����xt�vl޿+��;{_����}�^�4�ͬ����k�|�bL����^̏c%Ɠ �_�p�M��dH�l�HN�h���1��Z�r�%Q3t����E
�#��l�0�[1�܌iݨ����h�ַZ�ٸy���M/6>�,�|���e���`�!�l;?����D�ͩ�|�Nm��ėL/�2x�෌�Vg!��K�t�r�.t�oś;��r�[�1pn�uQ��zSD��}��'�$!���]K3�;/:�|���$,���&+�#文��N~��r�P��=M�	;F�҇#>ˤ��k\�Az�' yh�c%�' �qDkk���Vc��|@�Ǖ4�������΍�?�N4�귽��}�ߥ-� sǤ��i�F�����;mF�cdB7A(VW'O����.�{4�99q�s�|���a\����$������1�f&�����dJ���Ɠ�����.�������8~���O�L��R{�{�r�N�����)Y	�S08�����ڀ��[�i ��^5��7�����8W�-\���S`�A���zS���&��'<�܈S���@~�']F���5�--��s7c����j���hu�2`�����nu9Vdh��bt�g(Z9��A�R������uC�FĲl�@��fz�d�@WcC"�7�w��Z������Qt�ߍ�O>���_Ŵ����aw�P�`n1:/��+��2vdhpv���ELm��E�9�G=�}�~�^�n���I�}���K�����}v��#?����H&c�0џ���X�I�t����7
�������ݫ݃ྍ0�1��A��_qNS�bK7c*��`7N�1����q�N�vcS��߾���Fwk'��L���BҮ�^�/\��C^����`(�j��x��nrLǬn�d���e�i���JL��f#�e\�2���Ta��	7q	�DhF�=��W�"��*��M!�Z�n/~t6�_����&�J+�pJ���W��~
���N>�����T�T�(���,�ҹ&o60}u���F���')�@7�s��h"�-���Y��*s�줛����΍��P�B��NB?����!�<yⓓyݞ�����Sg#!;9�tY��0��㰂�t�gRP
��:�PFN40��Br��ǃ�GtS���(�MΙ�zx��a�FK&���'���'��;������u'��*�2=���3�AG��e���2Lfy��ʓx��O���׌l�l��G�~�1��/��
�����fW�5�Z͠.��h���tX�m���L6��g����_����to?ed.,/���I�s�f�w2����XZ]���2"^��������8��ە~�Gǚ�e������X�q-:�k�=�kDW�$�N<�"�%���.4�.ixQe���4.y�#O���u���S�B?���oEr�������lS�t2�	uJ���1w����x��;�9�Ş���?��O�����1T{9z�@�ȗ����}�(��<ގ�vc�:XT�5>Z->��܍����pk˟���$7�Yy��
�oA�G���J9�f�K�����vTmQih�.$mP4����V]Dꌬ#�R;����;���-JӒo���w�Ħ����/c�P�x7W��Y]*�s�,�DG�dE��A\,��t`���
?��5���Ntۭ�o� X^��|`Z?����v`i,��E9,]Xvt�4�J*�틕��V1��4�'9V&V}�8�r��m&r����ݻ+���h�ڵ�.O��c�0I�����N��2��'p1�0�+��3xb�U�v����>��0>k���0Y䟄�(�����=87����@'b�`����X�ûJ�Q��:l��鸓��`��9]�F�͠O�%Zi��ѝ�:�ߘ.yrШ��8_`���U J�@:iL6�۰�)�S���{�Dw��_jy�Ø�?�^���cŧ����Qt�Zs�����"*�gd�rǈ)ɱ����oNƺI�np$�ߑn�KCC�
�aU�j�ywJ�c�=�k:� ��%���)���� {�����w�l{����VW��'�����j�,��oum%�5��^���@��trp'�ټ�aKe--D��Z,�`�-�'
k37b|���	ɼ,S	�H9�~&��`.@V�+��'����׵���)h2N9ht���ؗ1�gz���wp,���������+���K1���gݘ��v��Q�[����PN�?ޑ��d#fz}�z�=�&�jn.���!q��2�w�����/]��k>{�	�Gqe��W��U������* ��s� Z���K��eǧ.�ٗ=�Ў��y)��+�۬�c�l&�gZ>�wZ�촌��z�{<^�ԺVe����$�,����	�kV8�������2��2�o=׾�����Z��g��̿�}��=V!7�%����e,{�Pr��
�"��4�����䛁�>���6-W�_�E�X�7e��:��HCk� ��K}�d�>�6L'���rI���ί�j9���(
ƐtG�t��C�=�s�����# :m��������CM̝������丣��O�k�Q�ɔ�Y�����d���JeRv\M�~uP=�4��D9X��Ay�h� �A��Yő�r a,49�g���el��1�،���(ِ}�����^4A3Q�t��(ݬ��i(�Ye�/�������'G�,�A�T� ���bC&8�u���_��!w�2����s��GA���bVe�������8���8��9-���|�{jq�G.Lu:���Ӥ98؋/>x?v���I��.ǩt7�2�܎�;�5!Ŝ�e%�tn6�k˱z�btX�a���r���H�Yk�0�_#��D8��6OȆ?#,;?�@ ��N�&�I��0�s��O�s;��������ū������W_�����QtC���ޓ�ȟt�s�^�W���h�-T�:we|݋�'2�2���bAmjz����?�#�Nۂ�F�I}��&���#?�#G\���'H�%>���O��v�q<8��ԉ��\�4��b�?��M��0P>�=����Y#z���6��� ce�����q�߆�l+��ޏ����������~ ��1� 5�Vq(�o=�?�)��!G�}^I��pfÐ*jp�t u���w��?��`<vB��^���"x���ˤXѡ=h����G�g{�ц1���o�XE��W��c�1��Y� Y�h�6=$w�w��a�-9??/��W��h�s����~�z�mpn�� ��F'|�����׮]��j���I�pF�G:/W�ܙO�t����sPJ?�r��;8�7S�o& �"O��$�4�4�cȡ�~���;q&{�{@d��}I9@ɨ���w�0D8�vcs#��>��5߉��&gb�24�UAg�z�B�,��x�G��Cs��`o$�)�IɁ���K��nؐ�1&���	�h�Ńdt��x�L]�[f������:��-N/פ�x;2*8�sF���ŋ2�4x�l�֧����Ǹ��ѓѱ&y珺��9��/��'������^t�����X�|!.]��V+�Ԇf��͠|�;��<[�(�
j�����.(ٌ3	�q]��|�"�t���SQ�=�QnE
/W1�Od �=�-��2fOg�T��i����X�aْQ�ږq�w�	�߹=�-�t���E{Fxu�&��`���mw׏�gd�1`x�iŢ����\tyA��ב�-Z�=rY�d��n�O�(�� �ע��I=T��+s��b����*<k>���/r����TmX�!!�?��zV���̣M�/�dՎ�C���ہp��۱��K������w�SK�J�+��1�O�L?0(l�AWqjj�1��W�,!��p^p��,�z�ߋxm}Ю����NG7��(�'�I<h&}�L�w�#D��e���|�r�}'��a�KV�,.�]2��L�^��Lkt�t��>>>�jF'����ʛ0����:8��V87���:��֖��h�yM��ޱ:gb� �;Y��O3�+_ӿ< �Sܤ�FWp�Χ�.5�y0Q8;2Q�A�ID�!F"�v���1i��!�+a��T�0�m#'�g�p7�S�M?�1x�qv�a�+�B�+�8�{G�<7�5mM�-6��>�	~`�:�&69�!eV)��|�c�M}�O@�ʫ8�7�N2)]�\�APP��u$�`c+�w�Ǟ���n���P�'m�P�K���S2[��ǣ�>����M�ܹ�}R!�a����{��86?�2�d��������;��kW/���J�{�8�����N�#�e��B@���1��F6�!1��U�;��!mR>�z�p��	�_�=��k�1����l'f�״��GO����G�h+�q��z^��+d�������S��A�`ۑv�����\3���6��r6��1G~�7�h���V��5iR;����bnm=��S�u-(�J���}n%��O�%nF%�u#<t6;#.��cF8�vZ�83/#��`Zg'�Q�ɟ�lJ6R������M�(�>���s�ԧ�e�N�qt�t��m=��,��B���"��ɏ�lI��,W]����]�aތ�p����Q�0(�}�dO
��0���l��]����7J�}ÊA��U1V�6c�Q}?��2���Qo	/<��~m��r��y�� iN8 W��qԯ����8����R����	����ꧭ1�+h�K2�=n;9`Lz�[e�:8��87������;x�	yttkkk��?�l�S�9��pV4��C�y1��#W�:��ŏ¯M����n;�$5:|�)&��d��v^͋&�fp�@W������ى�'�epbA�4�C2_~)ޟ��(>Ks���+����+1�8'cAw�2LO��脌S`��ѹ�������z��%�U���䄽\=��!|�(:!���'C�A�t7��o��gq́�4~@���d�-�~��f�d<?yU��,��������q���YZ�^o/���� �S�ƚT�fu�*8��0ζ�b��8���i���͔�7�$�Ho�z<~�0����ؐa���+20x�R��v��5�YЉ�T[�6Sm(�������(�Jr�<�=����&��w�c_�xgR�Q9'������M>]�ify>N[��x�������r���ޞ&(L�)�"����bye%�3'��L��zu;w�썓�{<��{2X�UGg�����`�Tۇg�ځ�=���nD���iY�SW�U�]�b�l(��Bm��fI|� �Xb�j
#�=�󋱸��9Z��X�M�Ջ��z�wt�<�%�7D�O� �?p33��'Å�у�K���O7~򃘾|9v��u��ҏ��Ϊ��uØ�ԥ�eջNӷ*�� /�ZoȘ��0xhk��8��֘��\�r���}T4�|*���G�h�?*W�mU�fH ��G���g��Qx�V�)#	$hT�Ic0YN�+id�I�Ϳqؐ�i�O::��8���,�/I����z�����[���w�9�s0��f{@~��_Ŷ���I����~&:���L���(:�S�Uͻ¤]�o<�1 ��2Ig� ����Z� �(5K�9�5�qZ��@��˟w�Y��9(_�T��PI�ߒ<�ͭ���wc������W>�{Y���������#Uv���Z�|�՘�~=��{q�՗b�ɢ'C�/�uVw��ɓ^=�.,����v��ǰh�����4�j��gs2�y�@?\=Y�o��d����Q�X�Q&�f�����D�2��~�y�=�v*�v�c����ܔq*#Lu:+���ߌ�矏+/�S��^�[�����`w?v����qLJ����'��b&�^t����Sy��ē�?�������� b��/]�Cm˛w��1	�^-���*��	D�b0(�ƥt�>A�!��4Y7�K3	�J�m5��A�<+�-��u�9>�C�=/��~/Ύ������_��_��|�I�ע��v�1���׾�x���y#�%;+2r{:�~0PK�nM��;��њ��ܽ�^��]�qM���/��2��u��T���zj�<~������չ���G��S�{�xv+�>p��io	��
�ޕ�x���s_˳�xi9^|�_��ʅ����[۱���G���+�p*�2��Э(�͊/�@[���+�C#�|%^�󿌛��qt.^W���d�������n�����ǥ���}�����4�)�c�c�)�u[��УuI{p-C���8cܤ=�7�ScW�Dw�ѣ�Q�b���C��`�����e�m]F�M���FS���v�4�,�Lj��gy9��_r�F���oߌ��2��?��D�c��+W��~��t����_�W<ߓq���_�Fؿ#�NS.=�O?�$>|������(�����NQ�g�E��R�I�9�?�=1(�?�U���8��Lؓ�(���.Ɛ�q;�~Z2�ѽw?�?�0��^�jbX�qqIGMteq���&x��x$�@v�Ѡ�	cn9��������7�w��{m�2�����g�B�3�=�z����Sa3���������NèР�I�:m�KNQ�'fAጝ$�\���,���nl߽'cl7��v��|Nm`I��s7lT��T�a�I���Fr�������U���V
ie�p��n/e������7L{6 f�x�wцČ�c	>5`{R�o�ǒ�'y�̲]):�F��ut#d��Ë|�O�s�F�R=���e�i�q"��=����Hanm�`��n�6o?�����qڡ&��+�~�>��Ft��?�q^�8�XՅ��dSq��2b���x��o��5�Q��\�Ӥ:�2�)��Iy�<W� �Jf�M�c��Ӕ=� �R�&j� �E����:�Ȯ3���������_���F�Q�C�MY�閏�����|;�վn�|·�v�����c�Ϊ���������7��Fi1Z���ݭO�*��  ��IDAT>�{��u<~��عs'N����ZXX�[ʧ��Q(Nf��G��l����1���+X����-�R7֛���iғ�)�p���������� D]����+����O�>v�j#I4H�p� ��'/.e��֤��qXi��f�@�E���k-�敕�mI��V^�7 ��L���_�Fؿ#���ar�H��믿�w�n,--��ƀ��^6�f� ��Xv�H
/��;Y��2�1�ҡ������U��4������4�3M��D7�9]�wvw7���:v>�8�2::�O$�����`�o�S�exr�pg'�?�y��j,:�az�[�2*ذ�[�5���G�CF�ś�c������ĉW>����\ޡ��+}Rđ��n�'P�G�7���G�3��`�W ��T%�����8��}`';2(dL�5�ax�V#�Z��%��Y����|~,���myp }i����G,���xa��O��ߋ8��S�/cD�
�*�h�/��⒙��;n���l[�\��]"s�9��９�*j�#0���N�L8�tdά�M�,���¼�ֈ�'�bwcU���:�~�ls�HUx�X�Y�a���vl�h=֍ �Ϧ���0�8��/]���4X^���o�ͷފ+��*ceN�R���z5Dy��]e��|#R����y ��қ�0���k��~�)e�m�/�*��֒�<�]��W'76��G��-���l��ڞi�E��h��,��o�s/�s�9�[2�$�@F]�K�]�~������ZWۘQ)���ۿ}?��/t�0�����[��������K���8T+�{�CE�Yu��<w�FT�I'��$��Ee��c<Ʋ|�M\��%͊#xYt3�$~��7�ɗ�]M�8�>��$�Sq�d�c��U��!)�3�Xе��[�@�'/��K?�:�h����1?�����MՆ�$��gy�-��upn��;:-K�\鐛���7�_l�?�'i�q|��	�պ���e�N寎Cg�?�6yMh:����"���O�h��W{���sэF0�ܦ���޽���8��E=��
�wcc h@������[\���vQ��d8:���_Ɨ��U|��_D�Ģ&��Yc2 ��<�;~|���}ּ=y67��_�a�S�<l�o �J��!����(���2�#硿��^�C���u�iY7�3���,H�rl�&�ue�n߻�|�F�)o0�"��a/��ёA6���d3��?&C�H�I��w����a��bo/�:2¦e��ʀJŨ�����Ps&mFr--��ڪ_)���@[+(,�mLyT����* g�(-u�ɴ�����+(���?��c�|lڟ�k��Ҟ��W��:��2%�Zm��{�����Q�ƚW�9�A?���gy8�� <82�2T���Lz�(��n���}W�kѹ|)�jc�ǧ~�����b�����B���b#Alt4n$oO�x]�5�A����U����|�b�I/mr�M
�M���^��{y3�g]�8siM��֏~dl�ޓ�~�a���|J���W_�W~�V\z������W����������oލ�緣�����4-��T}���zR�6:��97W�����I���6�j_@�"�Y���I��W�G��J<q�S�bl8�n�/�������o�]���5�'�4a��>��'t��V}F劯�B�G��K��8#|�T�$.�5�<�cQ��$݌i�Иp�f,��/����9|΍�G0���5Y��?W�>���t\���4ɰ�1T�b��A���l������q����M�o�e��A���5�dz�������tK˰G;�����bCn�������ϧ�A��
����a+18<���|���ƣ�ޏ�؊��m�L���G������܉�0fN��[\V}�4TpL��x˓����k0�#/ ٗ�9�=(��,��_�[��kp�@�t'O����QJ�՝'��`c#���j��ی���~d�{����	���%C�'�˘c�t^��˗���k~-��Ӭ �.��q�%�ɩ�|k�d(�)�O��t��A�+
,��M�I�ڞ*O~&1d����JC �Բ	��J���гb\��ze2A�y��h�?�iEJ���ffdx��i��sx��2���J�ϣ3>�C��`���UC�J�A2W5�f�q:���K���kq��o��_�N$W��aA��ޭ䇲�vJ�Pm��r�h��d�q��LJ�xt�zRw�]2��l]Э�O��*د�L��KOb �j�;���;�/��7߈���?���G������pg�+)e�E��/݊�\;~�U���ø��q������{1��m�_>��jn��A�������+�2�V.]���T,��I��\yc��I�se��̀�i`��=��[��;�/H��S@�i���ɗ���%����Q��S�K�nںM��o����9�_/���ς,���eJ��W�T���|!���u{1?7ﷆ�C<Pٟ�*��c���_�Fؿ#��3!��9K����a��ՉX�PǢ3��1���,�v�<���l'&� 畟���� a<F-Q@���N'훎��r���Մa����Gc���2 ��!�\=?S�o݊k��+K�q���?�$�a�>z�G�X�2P����>�t�d;lb��0�i�N���5N��೻�_�yl=�Tx%�0pũE��9D��mz ������:���3�&�H�`68�⌑���Dh��Á�<j;�]l_F���0Z��0o��X�ÇO�/=�(}�x�EHb\������t�R�lo���^��@�]��e%��D<�b�G�M�S�/��s7d��'s�		G:�^�Cn���j?4 6c\Y5���-|����+�ۡK��ʞQ��.H��✯��K22W��#�Ǳ��.k��\��Kw^!Pi�����(޶��y0}�j��a���?��!F�޸�~�v\���1�rtU��]58����?��1��&�n+%w�jG��{x��詇�\����+S�`�t��<�끌m�#G��7w����n�馤�K
��x��oyu��'���>�wY�2�۪�Όϔc����_�Ï>���oG����;���iVՂz�	�q:?_��2�d�ɨ_R�^X������l��ķ�){��lp�M�.�MR6��C;q��m�q5&��'�\�V�GYe��Mny�q�^�H(C��T����U~9׉h�W�(�M��/� �X��%h�9���8��S���^#x�f�H<������A�cM�Y&������&q��_�s#�P`�h������1�G}�|�i>~��=
�K��m���#���ЭA�:Pu���q@���$A�����@�O^s��:&&|�~�1Y&� �O$T�h�9�݋������=�g�^X���~+���9Mx�3��5���y�'�cJ�{���@e����~Li�� M)#:���K�"�������:����β&�Eݙ�֟��nYc��Z����@��\��Љe�|Ȃl�r�a�7�� Z�Sz�py���<qK�3s<�n{O���8v?��9w�jB3�A�hj�D��f���PLI��Ɠ�8o?vdl�J>�A�9_h�lG���՘�~%.~��x�G?p[��]��k�i'�F6-�Oݰ��v<	��N��R��䗓k�W����A�$@���<>mi�r~&e[<.,/ǵ�7�W^�ŕ�X���1̾�}��PXc%��Iلα�V;Z�}��)�P�'g3�kw�hi)��|��a-޸�f��j7-�=U���~N��nwm^����}���|��]e_6���KA�Py���>23��4�O�� �N^�򛘠�Wm�ǣ�[�K�*}iq%֗.�αn��������F{��A�������p��Sf%��ɴd������?ٌ���X����7(y3�Tr�����S�T��;���N�,��[T��G[}��sBSl��H<�1Ը�6#04��5�E>h=��[ap�?�F<�(�x�`�,�h�dEh�OZi�d:m~Ҡ��y|���D��D�g�YY�I\�B���Wq�O��ÿ�� �gl�v�����]Z�O���P�r�(Y
���?�o�s#�@�A� 3�d	w�ݍ>� ���s3gg�N��]�_��E]_���¿�#A��|�^���CW�'E��O9h�<~MJ���nV���������(N�b�3����W_��^~%Z2�zӳ��$�P��^?~�ƬM��#�*D���`��iG[����`g7��&���Ԭ&����??�sOX! ��ƞ1o�g����4<���g� A݅�#��rґ\�:�M�t�o�'9�B3�^%�����?��r]p�g��DyX�r�b�����8�QDOF\R3�沐WZ�����Ř�z9V��j����1��VR�0�~�V�9�7��)��G�E���ŋS�S~�MM���'�m+�:+W��O9&uVzfy���fM<���*�����e`�F���[�qtp��딐�5���H��d8����h�(���\y\-�W_{%^����_��Ǉ��5�u���T���;���b[�wVz\P}y�E���-�Q�d� ��^Sy���V��F��AZ�7�X��.s��aS�6	���L �OO�buEF6G���b\{��XXZ��;_��_�&�Ŝ�҂����>�q&l!�[���G��]�FY��qz��c�=e�����k =H/���D���a���M��>�U��jy�c�S d/�&Ǧ�㣶ִ'���8� U�@�qU�x|�V�B���?��$\G�
g����p��������Q�r��%�,Έ�SBT�e��c�&>!IߧM�x�����>:�6����o��1<>�1�a���A��s�'noo'~��_��:7�����38׀�Vy�'�!�N�����J�ul�fJx�GW£8����{�W<�AϏ5D>�<ɨ�g`DS?��Q�� :28��c����0N��}'o�u���yy%�28����ƣ8z�(e�q ���VI��<�b� �Fb���N{����8�ݠ��\+��o--�d)��j�`�q��w,��'_$�~t �VE� /���9:, ������|i�W�duc��UM^�9?R8��|c�0 %�ad�~�<"̠/:���iT�ٰ$?��2xt��?���X[��kq�ߋś7��td�0��mC�\�rz�Y�&TS9���h��Mˬ~ z�YW�O����G�@�$(C~��������v<����/bpx��w���� �)���h}=�?�|��vbjp]]�ϗ��R�ݸ7�v����
�rD#b��q�}�y<�������/[_~��u�<E�}��Is�K��3y�Ga���k�W�v��il�gҁ�<ҡ|Ƶjɧ4�Q��ވH�ә���_��ye-��ߋ�����˻�Q��G�el�N�->d�zg��ӂ�n�>�%�,���C<�o��c�CM���a��͸��q��ߍ�+>�>P��V�[�H�?�}%��e���L�ץ�*��GW�yg�>�YN���xCV��Ѓ��k��O���MM�M �	��0�n�c�o�,)�y�rF7qM�QA�7ڴ	�D:Ix�^�B�G�vZ����2�`����T�g���i87���2�pl��s�ۿ��x��q\�|ɝ�g�h ��E�'33�z�;�:2�_uX��)rpw"���ǂA^��O'n!��� iy��/���-�G.��D>ˍ�<���oFjP?�ڊ'_}�����̬4�z18:�5�1_\^�e;��'����q,��t�@w�2>�l�����&�Gc��N5A��m�Ƥ��$��k�j��`t��?f-�cnq�Qҏ�NO1�$�YG~Q��]��/Ô���Qs���LˁV��Z��Q]��f�B�2��>0Ħ:�X�t!.�z�g�����@����D{�m����?�]_�K�����ꀇ��$�ė�g��#��c�����O+o��l��8*�e���?���9��Ϳ~�p�pM�Kg@�G0�����)}�7�d�&lD�ͪ��eCQ���1o+��nǃ�>��w���a7�ȩtV{M�������x�;oĕ�W�h�0�2�0<\�"ٹ~Q؛��ߎ.������'��_���a���������N�����(̹n'�?m���W��	����ųC<9�9.9��=�l\ O�5�[�Q�AG��+ݝHF5�=y_��/����N��d��j�Wˇ��@���B;N�dLHǬЊ���LE��WVuc]��%��K/ĵ?�iܔ����q���V�!u2�b��4)������T��M�渤�.�@4�H*/��@iܨd݀�:6+����*'��(C�Q�-�5^�0�i?���/�����R6������<�)W�'���/4y����G�)��?y�\���s��pn��4rޡ&�����q��X��D� �������8��'�i�^P�G��L+�I`�o��^e�ݜ�$^3hx��D|�5�mp0X�G^V��2�����\;�}x��[q��Ӣ�����jbؕ����O���h�ۈ�1ƚ�ã��|\�v=�|�͸��rg{׫D�3o�������|{�4*�@�>���VcZ��	Ə�m�hR��0ar�x��}"(����M���P�br�^��PR܌.3���P5��)���¥��*Cl���(�}It8ߏ1N$���(��$��A�I����ϣ"&j��1���+?��7�ǵ�ss�?|�]��,\���O^�5���J��<��ő�?��̛0���>��5�G^�0���rY�du���?|
kN�N����v2���`~6V�����=�������ݻ���7����ze=^���?xKFG'6�=�{��{/��������8U�l�bo+⍣Q࡯>�q�Z^�9�i�0M�	Q't�n�x��%	�e��Q�kto$6.zQ�d�u#\�;E�0��I�e5�'%����>�4zw�4g����9�1y�������֖c��%ɴykyiY7J|����CM���fCy��Bp�J�����x��3ׯ����̢'�y��!0	�ג�`,;�tQ�U�b�=�3����ҸW�.����� ��.~n4�B\���?ʋ��A$I:����W֌��8����x(�f83e�����t��Pd�)[C&z�g��*���_�s#�X�Nܾ};>��S������@l�gHv �[^���#̫dB��FR����uO��M��* \�X��p��*ݨlwtᙫ�� ����%�����GI����a�i��������ǽؽ}'v�|��������Oc^�O���M��-,���j��GW��8�IF$Ol�)U��f�t��p�ʏf���j�����l.��_F�ؿ"�����P����PB��%�z��XϢ]:$\�4q	�{�Z��<��q�%��9m)�b/ĭ矏��;�~�^/7�� @�~�����8�4N���i��C:�c�1��D2�(�ɸ���Ɯ��Ź�i�fe�MלF�?8�Gw�Y�s���w���v"?�Hm����DZ�>�@{ ���ד��QĻ�Hs�l?��r��W�[�¬��I*qγ�����*���V����J3�kŋ?y;�����ի��d+>���|�P��@F�0�W����7�x%���q�����|����nlD�/G�D����n̫�x�+�<"W����h��6�:���	�O#�� ��m���F@�/(Ն�kG�L�H��&ul{R�Ǽ1z�flQS9k3�h�D��p�ȟ�C�G����_�^y)n��j\�v5n<wS�"��Me�B���ņ�;T��W����?����1}�z�ٽ��:cmmV��+��3)T 2�����7�<1ܾ�zսi7�A����R�c�3�ȋ��,���&S�|�7�'�J�8)Z��O�]�#��G<|����H���ЪvPO��#Q�r�ٓ���'�JɅ�|Xw.y��
/�,i�oH/�l��2��y87���@�u3տ�� �D>���ݎ�����)�{���0e,���}<��_�I�3 tx:]8��k:��z3���:[��(���S��cЪ��G�L�$��d0�#<�τ9�y1��P*���#Ȩ�����>-���E�-������Cws*ΆS�����
�q�;�7|��l�H�ٴ�ۗ�P2eTMk��FoFw�-�S<ob^�u+Ve��p8��d-�`01���J2�(����]�
��)��2Cr��Ifj�GD�K���%O��1P6��(�`��CHه�'�+M���6�x*>��1��(�߹[[�2 bAz�R[���36���Z\�s2..��P�✬)Y%g�N�������~�o�S뫮�%Q��ۊ�������G��>x7�ݏK�+����s됍Bp�Է�@&]	Ӝ<�4�A��ƨ䬛��/�s@���jYbQ�CHtx��U=�>P|gzq^FF+NSj'1����OW8l���ؾ�8��a|�����K_C�������b�/��u�������m2��m���Pbs��$��S��2��TO��x��y����Wb<��9����KW�v^�Ⱦ�>1:��c@&o^@�js����W��jw��8��Dm��XPd����q��G]�7ӎ�c��x�G?�W��_ƛ��׺iܺ{7�?�S��xeE�T��'�+ZS����/�K������+Wl��1��у�ٯ���Yy�Me�X?�<�"�
ye\���G9&��0��4.�!��1hp���B����-�'O�|@kl�g�q��'O�C�x�ld��8D�?iKŕQFY��1+�1Md�L��N�Fn��˗��F�0�'.��EF��<�( nJ��F2��7�����p��&�)���2vwv�׿�u��h��`̲�;��G�z[Ӊ�Q�:�ʀs'nh��8:Nŕ+��V��i�5x䥃Z ��>�xA���.<*���r�� �-6��ͱ�[yy�x�����{�G~�JcF�+CdVE���=�9�ş�@����cRʠ�eZiSþ&MԒa :�lN�d��q�7c��e���)���ۆ�Rmx_͙C>������%tA#W&JVM.U/�B����y��t4�̣�It��-���H5nhB���/�`wWz�+����.���|l<_���n܈�24Ei�����~;�b�|�x��ߏu��N1{܍��?�z����住b���c�p3��cV�-�;�15?G<�2�* �6��-,�J2�8���ʃ�ș} ���!'dV�y��~f�+��W��ʤ֙���q�v2߉��^�W��X�vIē���'�/c���'�����//?l=و�GO��ay��S��������o��-R��S�c��������4�Ⱦ"h�,��}��78L�uCS��nMr��8�q�4N����g�6�zX[\���E����>��ܵ��Ɵ�$���O�������>����?�ݏ>����+1-�_7Y�;2�j�o}7^�/��G1�6w$vN�ǹ��}Eʦ�Y�d<h������'^)'y��p3�p��F^As�HO�1�I "��ME*��?!�nA�:�w^�G�'y硭ӆ!����&O�-pi��/n�m����؄��7G�2^回��X>ݜu�h���C��|�{���I�s�v87���@۬�Yǣ�w�y'�ݻ�͑�2���r�:��/{�����f��c˗��:F�;��AO��Y� <J���\~��WwH����/\���k2�W��@C:��?cϛ�W�Fa���*}u}5V�V��W�<f��#ݰ2pD���s6�,�x��:-M�*���D���{Пm&$�a�qa1�5���N��~�S�W�^Ӥ��)��`w?�W�){�xs�s����2��d(ϕȆWY�r`��IØ��Ы�7�!�J	�;jb�}O+��������XlL� �gc�Ƶx�{oƋ����7��ۛ���sg��j|O�k�3n<=�7��{�ǝwލ��y?6��$nߍ�Ǜ1���^����<xe�ҵ˱7�c"L�Ȧ��(M�	�ՃQ�d\�A����t*�_�'�9H&c���z����f�cM�]x�f̭.���F�}y7�ޏ���h����IկW�D�{t�֩_�е���`c�M���1�n������VV��n��b�2��-�W6t-^S�t��i��^��$�!��NNH��I&YhO��P#84/����Se�mGtKxZ�����</���q��7����[��?�S����/�{�ﻞĂM�=֍OW�y[��ko/�����շߊ��8`�Ze�M����a�ҩW��.��B� ˕�E�ya��Г�TW�F[�-�q<�\尻!o~џ��Pʰ-�O��@�8;]�U֨=�S23�^ę�1ۆL�t�E��*ߠ0c��0���e���t#{�K~�q`uu�O;ȏ^���	 �Ҋ�s��pn�����>;3޼;���>�(�ܹ��˾��!���ø��A��3\HMu��u�󾭦\\�j��p���q'rT3X�&q��q�5a�еhxh������z�
��;r"��jJ�e8�]��	�-a��?��!�0p��?E� ��ǧ)�Ço�#�	�#/:�N�]T=M��J?�t)n��'��,�{.��T��I�3vE�'��e������&5�Q#�������ӕ��r�h��2�#��{����"h�'Gl,/�Wg�����kR�d������÷��K/Dw0�O�}?v�z ���bQ�����������û�ٯ~w�Nl��a�~r;��7�����b����^̢�s"]�A��9�j^)T��s� xG�(�����G�L�a2��L:x�V��Ky�+�\R�e�c��M�����t������G���gѻ� [;n�����j;�D�1�y��UV��Ay����U��I?�0EO�VWb���o��/����e�����NTN�.�(��
%� |���:��7����)�+�b K����1�Uw~)E��h�.���a�����7��ݿ�y��h]�������FO7H[j����W��_�K��/c��W�H���c>�^��`��+��+m�.��qIyF7(zH�3��m��/C�"�����㡝,�l�y� l� �1O�Si�5�}���Wmg$~���~�֘�e��<4��sZ����N�8��yV�h �Eٕ#���(�^��J+z��:�_x߆{	�F����6�pC�Ɠ'O�W���O!�^+��$��	�lee�w$���tO�%�g\:�S)	�Q�)"���{"S��jmN��h��SW�Ҧ'RL���*�]#|��	�Y��Ծd�n�}9����ڛߋ+�?3���ى���Mw��YoX�OD���+G7���d�� ݩ�C��B��CjB�������+������>����}_�LN�|�Y��]:��_�ъ��9�É�,��T��)��$zȘ�@�� ߏ�ɉ��.Yl�4iiJP��xh�X�Y�����o%�đԵ����2��>�\�Iww>�<��Y��a���2�g�G^\�"Z'�����������>�Ӎ�ht�Փ>���$/����w���Vr�رxa?ԥ��%�n$8��rg{¥XfD�?D�02z���z�}��'� e7Q2�w��LF���P��4�lHO��(��6c��<i~b/Sgfކ��u�j>y��a�2Ƽ�&�*�-���>�S�I=�������Ÿ���ͷߎ��C���0���__qp^}}�G�d��E�H����9��jp	�Fzv��%�����Μ��!+RR�L>�������������h?ފE�D�/c�/�]�j���2����ċ��Xy�..���@W�T��´%n��1�s�"ͻ�o�˃|)#�2Ӧ�_x������,F�Շ�ɴ\1rH�������Kҁv:3��LB���dcZc<�����?��>U��]Y&���\"�9:�^x��A�2�����J��� ��$_�$����N��΍�? �&���xi�L������{̫�����|$�:������qĽ�ʹ�r�F2�'��&:O]��~Mv��)a>��3יs<���7�b��gz �}9��knF�gcC�� G��K	���aA�8�y�}�ڕx����[�bp؍��M�Nq��o
j`������I�|�[~P��&����pЋ#�{����ċ����ђ���χ�>2:���:�nDb��̼����`� ���5u� :@VN;'�t���y��D�md���N�-��j*�%:�� `�kw{��g����+��ފ�/<o�>��o��G�����~/r�Lº)�-�G���֣G�s�a��bA���h�u���a2JOd��x�G�������B�J�Woܔ���S�։�H@76(pJ�]�V	�[a��7n����z渤�|M:��1��ù�8M��3�[��{zx����݇q&�����d��y8ӊ����wb~u9��Vb���h��M�'���J�.�A��Y(=Q?�
����K���~7~��h����X�r��C'����@�}E|��T;��D��@P:+�VF>�A'\��Ϛ�Ϊ�H�6�X��e�&�Zs�oJl�(ݿ}7�?�2N�~K�G�g^A=���1��̅�!��Gq��?���kq��0��ӳ����%+�禝�gD��j��Md�Q�'&dm�5�;iď�v����a� ��~�1'�v��,��S��rF��2���`#kį�'iC��.q�৴�l?慟���X�w������C�<f42��	���Z��<��E9ӓK}����v\�v�7�)_ҩk����/]���pn��A��UN>�����}�]wJ�����<n�Bj�F�)�y���7vu(�p��j��z����{��ɇ�iouN��gʯΉ�,�L�y�
�� ��#U[�(��AfM�'��4S�n��r^��W���?ڋ��51D����ۼ	�F.Y�c���r̭����J\��/�v��ݡ��[�q0����x�g?���W�Xt8�b�Aj?N�l���_Ƨ��El�g�=ˢ7-C��@^����9h�.�2��zk��g���h�Zf��7��7������@j�3a���N��_���R�>w-.�X�y%�2B?}������q�h��*���#E4�YB����Q7Z�����s�e���7���:j���aKf�q�������r,� �]�=ڞh�K&]1FY�#��Q\c�� CF�t���B|�=���	�Is;���Ldʫ/2�}�gϵ�v���cL7Eǽ��W�ʨ��v9�]��+����c��o�0�66��ʔ���/U�����`i1ڷnƵ?�q���?�Ko�sW���<�U6m��G.h��j~g�(��}�����o:��~G'����j�%�N)+P��ԙ&k��"��⼇�s܏���l���^D�9��$��Kq�'?�
����ԅ�4F�̴�d�o��W�0�O��n0-��أ�r�](�`N��!_��6�oR���F꒫�pdo�M��_�I#]��h<{e��K�^0���£ު���t����t�>�[e"?7Ĥ�w�Q<�N�lY<` 6�*����#I謰�QPeM³q%��sù�5~14t:ҧ�|����%_��0��v�u���k
���n�sx��l��z�@���L�P��0�m�G���+�y���L/�70�l�xq^郏P�����V�>����uS��A��tLwЋ㍍x,C��ǟG���qO��苎��l��y�U�����q��MM,���x���[�[���x��7���ߍ�lFmEKe�	�/����G���Gq�����>�1v'N{�������7�J�8V���-&��G͏@	^���Sd�dCYq�e�5a�tG��b� Ĝ�5��q��[����%;'�_x�z�]�(��$|�e<���8��^mFKz�O�L��� 2��d�����&�?�]���\�bn�pz����|lb_^�)�}��X�k�_���ue�#V�7�j�n�O���[;��O��?�O�Q��� �0�y�=H���0���ճ�ʇ�۱'5̿p#��z-^Q�x���bNF���^�om���N�� � >"=��>����&���~�}�?�F���E�R��[�>b���\{��,�s7��5OŁW��@�ԙ�! (|4:��D����c���a��
�fbia1��ww7���cC7,�l�r)^�뿌[2�V_}%ڗ/�I����v2+#��-��ц]�
`"X�(�V���@Nx��
dތ�l aڲ��� M�s��%�~W��!S��ť���@E�1^cp5@�i�k2O��r'�I\��d\��L���ҝ��	���b�)R�O�"\��pr3>�oJz��i�U��J�g�;��s#��28��}�޽��/��|t�4I�C�x1Hh�4[�	ʩ7}����.Q4x:������cEjt7&玩�:�����L����@��2�p9�:�骃�h4�������~�/S�e��ˢɛ���f�dRh�h?�~�E찡���1�������I��x���x����˯�*9O�Ƀ{���A��ǚTZѾ�^x1�jҸ���]����N���o�_�:�exm}�I������7�������__�L��ҭƧ<�I������.�Z|�� ��D ��֓��7�F�C]�	]�[u;�5�Q�&�iV��ֺ��8����(޹2¶?�2N�lE�5O%ϼ����D��#FK{n.ڝ�໠�����	y����LR��^�S/����b����b����1��M�g��d��v��_ʑL�[2�C��G>�<��~ꎺ�y��(��  ~'jO��N+.]��wO/.Ƶ7_������������?��ۻ��޳��/�K_G2���b��[������h߸]�Bюe~`�Iy2Z���d��%� a�c�7��xF^Ҭ�&��|�o�~eWC�O;�7���Od]�`J�:/��-�=����n<�� �:<���\�����O�!�Ώ%�$����B��	7R^e���8��Q��S'��c��7���5K�?�e%S���7@�!u8�Ytܞ����_78����gK?���q��͸��$�LK>*'�kS��	�#��3m��!{����<��<���&q�"ӈ�	 /����d���e�	����j�� ]�o�x&�+��a�F��'���G�����ߺs,�Β%�l�t�l�6f4"f�VCAW5��l�s �;=<&�ʸ~Ѡ�>�� ��/;�Dg��:�d\�x�<�7�).�[~� -;S9OJ$ ��i�-��H�q<FZ]]��9�x�҄���흘�0��J[�u#.��r|�G?�>�{_|w亇�6v�.]��/�Ͽ��x��W����_܎㯾����6��� �����8�܊N��G�1��yOo.�.G�3�ɴ1�P;��P��,�r��HWT�@2���A�@�Ə��GW������=j�gBe���w�b�����}Ô&�YYQ�;m�Io�c:��ŧ�/\��2b�.]�~������e�.nDR��Pg�e���k�ĕ� ֿ�ftn>ǳ�į	a��dQz@��� g��oL�Ð��'�����n<F��@��>8�Y_�>W����/���/���qee97���e<��v�r��~�v�8nXU��N]���x�?�u\���c��%�='��{��Y*1�)�F���#_��X`��9t�,HWx�嗗��A�����,�ZA�q0BгxP����F��P��X�;�Q��g�YJ�5c#�xe!�}��x��~��nI��j*�	Y�3T�AA9�{�m [��$�oyh���_#j�jY]SN�������[�Mm��F�yC�F��FRir���y�ׂ��J��W�q&��O׃���I�I��-��E߬��0��&�r�Ccp_|���c�+y������{�R�J���l �ٲ������������/�������: }V�Ũ���h��ֈ}g�N�$�	�G`c|��q �c�c@�]h�iG��tp�<8����<�0�wPe%����8ʩ��Y���`�1�a^wc�不V���M���K�6�敲��DƑ����+kq����o���B|������`{S#wy3�YZ���Wc��?z۾�0>���;��u���:�7�uԋ3/��ik2ф�|G��8�v������^^�a�c�"F_)O�/r��F�U���qM8�<I�1.�^֣&�)�O��:'V�j�cuY��b�$z�8�ۋ��N����zB1���Ǻ�\���^�e��l{{�q�>��1S�&�Y�q$FT7��/��[ߑ�v\����s�zgd�ql<�)�� ��d�[������J�I>�R3c(yG+Gr���4�CnP*o�N˨�SN.�?�_x��9����R��(�)���$�~�Q�����ػ}/�6vm�qH+�YAۓ~�`���d�����ŅW_���\l� =9����vt��R>��*��j����9�]p���c��F��!�8������i�?��Y.�A��:�
p�v�X�c���Ho>�N8���}h�yQ���q�%�7n���B�e����W���mWep� �|�����Tc��y���Yё�Z��7`��F�M�����re�~
__ݞ���J2�ܤ��$���nӀ�(# � ��1�9�*}���8Eer����P�YOؤc8��UA`\󓴀2NI � ʅyq����E�_�G����;��s#�M[�q��r_��ʊ?'�GJ܁����n�ƜW��8�� �F��;�0&.�: i�p����aj�����:�~����J7�W��<�p��! 3��9�ϻ\\)�V�J��Xx3��&X�1� >��᢭�vƁ�;2�n�x�//�����m�����{/��Æ�CW=M�����d3��y�޹'�7����A7{{����1kR� ˡ��Sz��e��Ȩ��2w��֥X�n򏀅�� \�R9�/t�rJ�JRb3q:.uW��	&��0?V4�oD��c@�cE���Ϸ���Tr�v��lq5�_� 9@ƿ�o~'^�ޛq���X]Z�Ml�}�Q��lřn�1<dL�4{k ,/�c��~��x�?�u���Z�I�)�eggX���l�n�n� {)'+9��āNr%�}(l�fÙ38b���Dn�m\^�0:`@X��Q��E�W%�@�
��O��nW���rt:��/�������bF���@�R����T9�N+��$������~����)�!��=��|���iK�e�[�|'uF:�����f�mG�R� ?�(5d<�f��O�YFpWq���Ġ�gD��C@��h��(�E��hK&	�Ǉ�7��]����hi��?�~�v��VB����j#L�vI[���[���f�D4�"����\��� ����ź�vj;FxıW��K��F�O̊an�M�k��rp��a�&4m�D;�� �DM���m��YO�]����t�ǃ�o��Z�"eM:V�l<	��֑ʔ% ψgɿ��>q } |��q���F\�r�q�������8�@P��z	�[��s�����ofD����O�7!9�����@��:��|��NX���8tM[$���p��;��|��MB�/ �� U��� ��|�b@�|?�L�ٹs+#���<�?;�'nEd���AE�2��Z�鬌�{����|���?|��8�܎�?�O��������m��t(r�ua�aOF��
M�h���o�1𨊏d�Ȏ�9�Iӄ���kOGwm!.|��X��_��w��/_N#Cu����O��ё����?5I�FX���@j�t���<My1�"G;Ԡ��1p|�_݉�|��Do?�߼7����˱��q|�7����Ν;���'�y`k�������&ܵ���B��h�ņ7����:10�5NU�ֳ'�c��@[����Ɛ#m��+o�#n��IM;+B�%~��*�Q� a�y5�#������}ݿ����'���Q/E�xS����Nbpq5�_}1.���������1s�wH� x�~]�4������u��A�}39O���+���]~� ����uO�ބK_�xJ�8�Z���d̛HA�5�t�ڬe�I��
��s�ʤ&`lP��,����*S`�F��9��*��Zd���0�d�o!��U��?*,œX.�'�x�@z�U���k���yO�|���8����_�zoڑ�$�W��3�x�/�A[�8���|Q/�tț7�(���|v�[��[�n5���p�m���o������O΍��N@��8t$�\�/����I%CV5�A�S�ӹp�E���T^�8w�V|5r�/�D�/��ř��2���,��fL`pj�����V�Q2=�Q9��s�h��;sE�!��ߋa�(�V5�l~�I���_��_�í-�N}���~5���OLN�
��d���C��Ū��Y*�p�'�����߉�?�����_�v=��h��c��rXxn�\�9\�
Jv_��9&�F�i�2�o�T�iJH4�0�8�ã8�ߏG��ݽ�t�B�|����Q�)c��_�2�����mGq�=��Z�W�������b�1>��x-ڗ.�0Q��,4����"6{bV{�O����ū�DPW�����aY7�g���SZ�*��h���~��o��|�� ү������o����)���q���X싦2�η��8�o����q�{ߍ��Hmd �}��e�+W�2�甅�6RF� ?2ٗ�����Q�uW�k��/aڅW��?҇q���9�T��(����0"��c��c�&�ęo9���Yf����W��l*We����I���G�2R�3���Uv��� g�Yr�O�eY2��5�f:y�K��(������� ����%�*S�O�44Ս'Y�]��>�@�˼}A.�������a�X��>�^�$��[ԕG��?�яbnn�2�.X5�r�HCǴ9tu�����;�ND�으a������!�c:e<8��F�F-������V~������3gǳ󠒎4@!_�3~4�iu%�d��NE���_��>��k�� ̸�\�פ!���?�r�*xy�֠p��[_܎��'��k��h ����c�b@l��fZr��0����	����`�<����P��k`��u3n���x��~_}=��l,0��~Ŧ:�'A�My���H&��! �[qH�1T>hp�W�.'
e�z���W8�,]���cma!6�޳v��������O{īA�3��H������ߎ����ƫ1�J�P�Ô�L�pD�!;�^��=S�6�& �D=�~̻��۳@�������$��ǳ`�M<�����N��l��l��x�p#�G�h�����7c��W����8.��Z,\��|�~�}&^)��/?�����2��Ϝ�͕�I:�k��|��)1��r�����=YG��?�]�'Ӝї��3�W�'>Q��T��o��Z8�E�h'~A��a;Γ�d8!=�cB��8��s@�K��:ɽc9�B��f��:i���EK���t����&�� y5m�c<��䟯U�To~�:(�(��U��d() ����S�C;�����+��������b,-.�p��`^���FؿTǜ��؀��'����}~n�{Th���|�~��N�el��Vu
\NT�]e��q��@cPp2ﷁ��g~����2��6Ptj©N�Wd�q�d��]������@ʝy�/��.Χ�3hh����ã��ɧq�����믣�p��:&=�Mw:q�)�w:ۊ����,�[���/#l�m��>o?*8XZ��o�p������­�^Z�fu�I �L�o\' i��S=�a�'�t���9!�C�Է]&�ϕ�X ��9��Ҁr�{O~N8���=������ч����nt��=:
��q���Px�]��͸�g?�+?�~���r���DWt����f1�a�d���W&��m"O���L�Յ�ViU�e� \Gyu)��'�x�7�
;������Z�����s�fڱ�{�6����q������ .~��8�s<|=a(^����M[P��u�_����r����1����v����u$�(N�M�x"��o�f|��@��r=	̏ W_��J����W�2���h�8ؙoҟ��6t�\_�rs�ɱ ��O�]�^�+�lT��F^9�����C�ɤ�����k,;���,#��@�J����ډ_}"�V�ɇ��D�/��HsM��o��x�&N89'�1
Y���h����2ƍ7�g�_�s`>W�?ek�~�P��Zڵ���,�����w�˺��F�:5À���C~:�hT#'�j:����gp >��
LWP�� 8���']�K'��� ۔�k%8�~�$G�HUPPB����Z]�h!�q�''<�<�EM��uEpVFUgm%f�d�G�q4{���+���_�n=�_z9�kb�p�7�#���L}�?���N�W]�ﵗ���~W��V,��b�򚌛���q'��@yGz*��g�-��9��$.�:��h�aS�
�'	w��_�<�|���@����h�}���]���^�gg�'C�?��Ͽ~��������/�`a1�Tֱ�e��t����f�<1�ã߂xe�I3�
���䔋�&��P�rd���7m���	,�P��3�~�]>����)�X�ޗ��W��S<�~�v\��[q����ꋪ��y�=�baH�����Y�I��9�l$8�8�q�f��%��I��
��۴�K:j���7e;����9�QN��66.+���\]ӟ��ʓr��FN ė+��t��+�fI;!�(�@�1�.�����:S۱S!��G�%_�dy��K�<Ĺ9�&Ꚑt��Zx���ʅoꘕ8�pU:�:�z)M:�cuS0J#,����E?�=��@�5�$��>�ۑ|�lo�������x�渌?U8_	�}C5��J���3�q�����9VWW���ڞ0�хO��fuukw�lN&l�k�iܾ[�U�z
����	������	��=a���[T�C΂�0���rU`c����V>V��)B���H�o�U�����̬Bq��)%����BHӱ���ۛ����_Z����X�v%V�_��7o�-�7�GGw~���8�ڊ��_�m�r(B�pO��ˋѺuӏ�n��Oc���Q)z⛏���֑���D�R>2�<�5x)�XG��܄�ڳ��3���<žY��(�����c�l|o�;1��X���Ǜ1�ًӃ���]��b��:���+��_�U\�ɏ%�s�?�3?*�O���w�E�vJK�&��M�Ot���э��|�Ǉd��T;+���*�q�QM���|i���hOb�'���+�
�%���B̯����˱p�R�]\����4��	_ƨ�N�� *�ˏ��4�4�Ӝ�D�N��7t �Q��x��G�ɉ���y��Y�W�b�&~�%�g��&yO���lI��8�2��eJ\��(�)W���j,�J� �����6R�H���>I�0z���I���S���LZFs\��1�0�˼��ٔO?�p>R����8�<����Yv��T\�Y镆��,?�.|��(�7��_���}ǜ�~\�|�y3=s�.(>�*�O�7����AK�*;2;j�����{�N\�r��s�ꮕ�X���R���0qx�䷞���VW�d�Nv<��'���J&��fu�������M��+��t�G��+���HO^�) � �f�����)Ќ��D��l�d�r��q|���/��8�َ��Z\�v-.�_��kc�G���*�|��8x�$��ݘ� 7���?�<n,-��k/��}?.���X|�9A N�5���k��]��s�#V�!yՉ']!X6�X=�g]����M4l�F�GT�#�ep�.�r��+`��D!˂����3³2��ލ�_�_��?F��;bJ��.$��_.^�ٟ��7ߌ��KqҒ�j�l&O�0�t���4�o!T��J�~��mY���t���5�n���<�gf�n�	��A���4\��15��O���<��̴T�EW�� 䦥Wȁ���uR�J��kG�?������Lʑ�<�A\��|�a��4�F��V��mS�vqc�b�.uU�)�<a'��gq����'�_����|�dZ�Q6q6��q|�#obN��0L�/�4�B�_Jv��7I����&�%��1B�:/<]|ʧ���e�V�g��I�(���!��S�|5�!�CSe�;Q[˽����n09�6h���7eɯ@����u_n�|V�(�.j���?���w�+ݵ|tF���懂o��O �W�~�ྖٍX��c"h�|�׿�U\���C��9�����ݘ�}\5�:�d�-y��e@�
�٩�n��<�g]�be箰�	��G	��F�r:�0��IG�
�hd٤r4���L�B<=�ֽfz��T�[�D���M��ҍ��6�o��ݺK����ۋ_|_~�a<��eLSo"���Oy��Y�c�y���o�/�����ގ��+�c@�������Y���-�x�+����#��. ����1�ĕ2O�qWM>t&g�K��+z��o7�eL����0onFW�֜�՗^�~�����[ѹv5�4���hKt9�}A�t��+V��q��YW�G�Ea�Ez
�>�^���� �w��#n2?za!W��:Z]�s���R�Ǿ���+�)-{FV׌�@f��uL�u��e�Uz�7KO���$��#@��U�2������q~��3�V�@�+>����ꓲ�'8��U�zѪ�8_�g<���8�SGI���f��y���q�����ax^�D
m(� ٮƼ"#0i�@��DIY�,��@� ��Sf�����
�A* ���.0�^�5�P��C�?Y.��>���p�4�N[�F%	𓺀,�|U�s�k��_�ׂI�������Lq6 �Tף�����ފ��������n�0c/�:��ec�C��J����1��DC����;F�Ɉ��4�'��$γP�\�w�&���	��YeeG��O�ku��� ���r�}��v8F{\��� ��TS+`^�{�����dHp�(GW�� Ά�X'[;q�w�!��=��?�����t=�¥�nve5��.G��U�p�;�F�ҥ��̭��L��zL�ݿ�ߥó8%�����7Rq�.��v���W�B�Վ��4m@��Ojq�m��<�����^<��Ӹ��w���0.]�/��f\z�8���cY<�%߬���.�C~{"�?�m����p%=�6����֛�+��3���x�\*�0��+G�~<�4��H����F�OE�d���I>$�V[i����x&>]4�MZ�8꤀2�$�Ց��}�Ӥ1���I�����'�?.ҕI�;ҋ��1h��w9�6�;�k�������9��^���ʠW��9y7!���q��������W*Oa���l� �1� �V�
���*L9��)+�ن
�΄� oi�$�f�e]rE��W�mȘ~�6�����cp�;�*�@]�XJ�|�����?y��p�(�&��ғ4e��֯ނ�"#��&?�\C��,���*ZU��2�����
�F��8���K���]���~����œ��q�����'��Z�d'��Da�	�/�tE�	T㭻�D���g�M:��)g2���w��'M� ��)<������M�"�<to�m��ӹ�Wy�oy�0�fb���O�lH7%g,���h�qi&!�0�����vl޾��[}|�ݾ�d0�Km��N�H���eo>������/��7�li1��"��:��OXI:�d��-��b�{�p����A����!O����?�gd�
�&:b����i-�>sr���H�
���t�Li�3#cc�׏��O�pg'ں�X{�z�./��������#	�&�lʥ9���j�x�A][����~Q��A��	�n�/�4r��Qv��?K��yk�U�UL�9��%o��З���ǥ��ԭ�p�e �(�*�u�+|�>��ʮ��Fg�GuUƗUՐr_��u���J��R�i8_���|�3C��aJ�@Y��,�f2y��m3h�M��w�v�Ve�����є��Fej�d�fuڬ��8E�!xĕ1E�,b\r�OC�����_�H�����I��@(���;� ���}x�.7|��n5�c��"�<"��4x���G���C��?�&%��1C�#�]6(�x�@,//ū��&ܖʪ��2@�2I���O΍��'�I�l�\����.>���x�������1U��f��d��=��/A������t�jĕF�:0���F�mP��<EH��|T9���+�k�K�[{���/P�HX12�/(�I`����Q��:b�9��� ��WAƋB13��������&��2��ߍu��{�$κ�>��G�!����K/�͟�,�|����v)���3�
ȩ&a�jY4Xa�T5�9߭6�VX:&��#��:#>�����OB���3a?"xuJ��Þʧ}0h��t�y%��p��=�9<F[z��A�V�#�V|����z���4o�'�؟�a<��F�/�s���t��6U�n���A�V��į�T���%��l�'��_(�y+nt���hҡn؋h�^�;�~.t����ɲ�O���ơN��0�"�~��|n'r����	��V\8�b��b�j�Gxiʐ�tKS.��A"^�I�m�)Hy1�(�7�1j��)��f��݂4���H�6�'��1@{"\��h���v�������b.����+��A��J7	l�`u*�!�"�>
rW;�@T�tQ}��We��d�������ÓP�(�j�@�d���"`>���O@��s'��nXeT׸��Mu!�?-ߞ�z|饗�K*�h�뀼���O�4��� �<BRc��Bق#�޹��y\�zՃSJ8w>~�6!�dGs|u��ѱ�t�LKti��d� ��:�;��L]��7tk  H�Spe�#�e#�3��;*�� �7�C3���*\�쟠=��3?haF@O�r��d�qM0��g�r�|�r�r\�v5��~t��c��Fz}��#���B�ݸ7�������W\��c����ei�cKu�dG9�D��h5��'2��ПB�c���O��/�uY��+���"�6Su�Mה�A�.�:U�U~a���	֯��#��r#�!>�}]�ߏ��b�J�>oM�o&2a�G}W�]��WA�}������%���e�u���
*��ă_t�F��̛��p�*8�j&�]g�u����0��Oa@�H��h%d٤%ג�t�xR��ґ�mD|�T�e��)L���R�0����?��i��x��
ߍ�0�k���v�_����u�/V4+7�%�h�
��"�p�5!� �>tM�L�Wry|�����,W����FBY:*�}r�hi��M{5�,� y�_d��p���Ǽ& /y��5���c��i(\�ڰ���o�����a�ǚ-ѥ~	���&L֣��|e���r�BY����/�&ɀ�?y���a$+�nj|���,˅����J�?�*&�ݷ@!�c�q�&�%������=aG��.�݆4bƢ�8ٍ�a� j�*�R̸��W+M5X�j��S>�$�& \�f�+���d��@5�s���c���ɕ�ʤQ�"kRt~25e�_^�/r���JK�E�����C�'�?��6<�������]��ۿ�量b^w�<*>��~��X���q��ߏ�矏������Ђg�/�)�t�b�ulB�� �<��xZ�� e����/y ��-���eA����Kw�~W�*��\q���N�Q�9�g�I(<?^����o�)��I�z�6}O�Y��O���I9I��T�d|N��ϊi�ŵ�\+ŕ�4��T�	��u��n�+|��e�YA��3��5'2P�e��~.\&��3�8`���1oL��sv�.�(��˥���t.*�SqWap��B��?㓆y�8�[��'Їߊ��=<F>e�I�/�&dn)~�1���L�}��M�g:Ӻy��x�~0Δ9�.6<e;��+��_�:���|&�O˄����e�/�I�:��y, (��tT�Á�I�yË�&�04�o�<��$���*�V��%���2n��ƛjs|��i���,Ty\�d�S�q-��;�C�2�����n����n\5Ix�T�́6t6�qU��(W�.����"?��!<a��#n�0�oʨrH/Wŏ4�N>6��f�V�PWp �7n~�lhQi.��ɼ�~7<U:PW ��� d��L���q��7b��q���8^��/����_�w����+/���h@/������ZȲ�<�'���T��� �W}X�
��r<F�2�#�e�Jz�&����QJ����t�md����/�g�ڇ�Q8�gӿ�?�[��d���#O�����Q��gp̭�`VYM��t��|eL�|��T<@>�%ǳ0�_:)��.�gqU��g��WP��_��!/H	}]�S����G�Y���p��%�'閟�r�W���*��$a5����;��$4��k�
%m�\��\����S�Ø��Plsԉ�����x���-�*uYu�>8���n������93㲕�6�csoP��q�m���ӈ���L��ȸ�q�𔢎��'iٞ�_u�ڄ�"<��R�3�<"T��:�d��j��m��;��8���ɶX�����
��7�Fꐛ��m���`TvѬ��H���)������h�����_|����~5D�����A�г�T$�ku�
��]�<I�T8�{k�#�`&��I�&ZEW�-�ܺέ���t�ʰ(��¯	p���p�o_��%�M�!���RA�|��D��XPt��bQ�����t�⠯Dto>���^�������7��ny#���2�gY��L��pƋ�q'�8G5����)t�t���T�$j�)�����4�K��I���-@ZMF���˹-	J���>p�䳍o��7� �FH��\1.����)'�(�>�|6f�x��M7��ϧ�5a�]����g\�r-}�����'�f<"�0~�y\U�rO����^	B�(0���g������L[^�O鵈L eN��+��i8���y��oF��tNo�׉F=�E�ݱ!6�wc�3��O��_��>����tn�z>�4��.�%D���g'�Y>�V�N�����4d�7㉛�whe=gZ������_(~��|XC�|
�+f�^mH	���&PyL�)cī~�|W������ӕ�E_Ѝ,~hM���`��?%87��+�[�Q�� ���F����_~�����L�٨=�)��Y��D�&-�|��0� @پ�h�p���U�w�p<~�5�9�%}z���� ����>NHv�1]�P4�D��iܹ�D��?��&'\ 9β��,����p�xq��xzpɁ"�
?0Ԡ��,��ƥk7bn�BL��Ǖ�^�+o~'�o^�n{6�\$oK�4`��1蔡PB�R�SY������y������zD��y�K9���
;?xd��p�ɛ|�n7*W@xR��Kڤ+��QxM��OB�5���qM��Ys��T@ч�d<�t(��F��.?�|��\P�&��/Y'�>�SnRG7��2�֒�4��U�zv��#{�0N��_n.0ZX-�Uad�5�IOjÖUtre(������H�� �7���tġ'2.�+�zn��k�G������d:�-�f�#��x�ڙ���G��·��'��懟����bmm-�{하^Y��` k��NH�$o�ZfN���:>�FS�?y�t�M��$t�Sc����z��Z�!b>H�O��'�4�+.�	Oi���) �^�PdƑO<՘�D�ڇ�m�?y0�X��,L^�X�XZc�����mP��u�S�q8��j���������~����ύ|}}-si�?����o���F��������L��xE@���4G�Sa�OB��
�y�w�-�v5�����F+Я�E����x?�á�K�?��+q��r2�;<~M��R����Hh��;��^�_K�`э���~w:q�o������/b��W�?7=ՠ�`$B�_S���3rЗ@�١_<Ȫ��o������KjɅ��.��u��op�l38&�w��Y���[�bLg\�E��d{���|�����K���	8�]�ʷ�e5M�J�u�0��$�O�ʷ��rU|QV� ��	e��\��&�)�p��j��7A�z��P����Y�pÈ�,�םH�C��tI~>Fϩ�*�k��R�'��ن��M׌cE�Ʉ�[�'��xҞvi��տ�A�� �OW�	~p�g|��.��L+f��+������ ��<��G��dg/��ߏ㣃�i�h�����*�t�>���83S�r%�7�9��r�'�J��{%[�ʽo��h�W��}BN�|��U��:FOI��O7��Gq����%�8�,��Mܨ���:[-0p�|�ȶ�/a#��������5}�*x��0`����}76�6�u4���qR�;���HG�?�!�'ΉJ0�Ə3�������|9͝��7y��չ�<�g� �I�t.[W��p>\�3/�0��>�11)��`¯�F� �Ow����1Qf�(� 
%���`���jk 捿C��elM������$��QՄ>r �FFW�c�2�_��5CsQ�@������[� ��m�/�姮H��A0��o\~�z�A7�?i8���Wy�J#�S
� ��7�~'�G~�X��ҁ����ⱜ8�U���b���}C ��	��x܇'~�W�?g2C�����M�h�e�d���%?����/鈮9deLc�⸂�M�]�o^��'җ�G�ӷ=<�%թ~*���R$��፸�M*)[�}Ғo���i���y��ϸL�\'����gO%c�L�@�Q�h�z⋣c�/�ҥ�z�b�O��[������#o��K&���ѹe�o��ה�ܒ=�)7W��� qȝ������K�]�/���PB��̯��y&q�j6}Ԯ)p>��+/�TmH���CO�sp�xxx��%Ty���K��T`��s�W��B'��q����_ŧ�~:2�h��&N�w@un��Γ0�ؓ�h�]��>ˣ��@1n�9x�廓�A�ɰiW� �h'r��\�]t<�L�7��o@)O]�/�ſ'P�E�L�Д�ō����T��P	��pY?Y>�#�*�I��qJ�w"98�u ?b�ҕ��ԁ��rCA�X� �ʜ���S���O�2�A�|�U*�Un"�N\�Yf�QJ�f����?�
���]��)(~��T��t�Õ_�^ꪑ�8��� ቲ�7c9�Ɓ�\�˔�=�r� �-RvCk�W��䇷j���:n�p��4����:�RR�h1N�J��Dy6N�`^k�t���N���y�
s�+D�H\d��4��~�8�3���p�
c�<�A�>'M�z����z��Ue��~���#6�HFO�!�72�#9ň�2ڈO�΢I���0�z=����#�3�����=>7{2ӊ��K����՗_��/<s��c�@��ޞW��C�"#F�4ﾗE�GS�6��x�NU�\��p�y1!�.��>Pq�#H��EJF�&C�� ����&H��F�n�X �x�_����,�?V�T·��Yo�sɒ���������'Ir$�� ��irV�5'�=3;o�ޓ�/�Ȼ��#o�vv�g�T'Y�yfp�4"������gvu��o�խ�
��B���`#:@�!O
&�'��-�Xs��)�pT�N��}���队�cL��3�� 'xL�6���Fvs.��F�<p+8]'��\x
��� c&��:N���s����`�r}�N�\�$�OY:#@Z�}�&rّX�b1��������K�/ë���
	UG���Y���^��ix��) �kV�A����T�5G�d=ԃ�Uk�)(��eB���0�e�t5���\p��=;�n#�<S�>Ǧ	�{���jW�&�%�]�G��+��*-�؂sH�G�"?��O9$QR9�1!zeV 	�1q���, ��N�ʣ[�{�s^�>)ɘ�a&��S<9����	-�>q�	���&��C������|���s�q4=�>���Ύ�y�� �m�c�5sm��N����|�kV���ӡ�s����<��j��n�6�q��^y└r���2�P,qY���8�O�`_�v7|�ˊ'O3��x͝bY�̇�O�Iv�0���cnm3.��~������ߌ��B�zʤ}�]Y��v`��}��� �XȈM��ǔ�4=��-����sR�#h��o��	 ����6�N/���F��x��/�I~�^�i��3�&�@QΡ�������)�i��՜�1^�D��`�N��Z�+��}�����2#��+����m<x�0VWdt���@���@Yvs^i��uNѼ������A:)��&�� #z6����&��ͳΫ~�jRz�s���U�W�a��.��ଉI��#\~��&�����M�?�t~Jf`�������	}��m4az�I�\m{2P	�|��a�C_��?dBd�|�� .e�����N�3	v^�:,Aq���	������i��$Wb(K{T� 瓀,���
��`�&��*;���N�O�.T*�}b;�D�ɟ:Lm�Fвav����Ϡ2����Oɥ3&�񊆱F��9�H�f�fu �I����#����h���$�~NX�ґzlO�q��e�cO]��I~��/�E�����0�{�q�����rHV|+OTU��¦XRe9�����Y�v?��,yK���㫎W���l���*ol �A�ӱ�<3�rv�3G<u��ջ(���8�u�v'��=�Y0I7�'z(*�=;�%E�;����_�¥�q���c8j�=UdjVc�<8nSR?r���}#��A�m)#��2r�\�*�Qڎc��э��I� ��-:��4pHi�I~(�����zy7&�l��R�	U�$`����7��/�Hf�. �r*I#��t:Ν;���˶;��=	�Q��[��;a^U̫&�2��o��/>��oCr��q�Nl��_]����a���D�G��@2��q�'�u�CӝK?.R}��3�s%�r����c�9�kũ�+3`T����Ov@�(G�:��M:a���8˼1�zHW�M�S�:$o�a��������|��5��nhԻËo���2�X�x�E��&G��&���W+[�>��2���FW�Wtg�QX�F�5��U�xv���#6K�����N�>����#C��Ԅ�KH<l�e璕V��,�5�t���A��_?�Y�E���j'ˮ�$G���0nC��T0rʛ4�2��`w�Y ��|Ɂ
�N��_vB~	з�'��Iݕs��кK}f��r��[1x�,�w�c��E�t�����~��+�q���>���b(��CS*L{�2��\x��#���`BG��1�ld������[��+ ?�X�T{Q����/N�cF2������{����8:>�sr���oze#�j
��M[��e��I?�ں�P����=�~��Q�_ϙ�3�ن �)�!��<�ݐ��3����H��ݹT�?l��/�����W;�L��V�$�β,���8)�ǸpA�@�dL��s��3��[uA'��K*x�q�e�~��_^��)��«1�o��E�����aoo/>��ct����8Ӹ&C��ǯ:i
��{���Y3��c��Q�NT8��q)W|��֔%�����8����7u��S^Q���M�SY���5	>տg��WӒf�u�Ш���}��é��� ?,�0��X��	*')2������*�����M�x%k�c�W�h�o��p%�%���h�Q�rʊ��7+9`fz��W������'s�~?w?�L����礊L����N��4*�q2d_�\�<��v0d�U���ܣ���e8��� xb����2�x���
��ҷq�c��P���I����S�o\~ds��!ndz�L�q�&����������@��{ѓ�����0��0���6���D��8?���܌��N��cni1Z��Ҿ����JY�8����U�j邼���|dz���OQh��+�P-tTv�D�vْ��Z�cANR�ν�q������>��m9�beIr-����P�Է[g
�ɇ���]��37����\W�{"���E�I��/������p:����X@�b����XgՎ�q*�D֑�:*�J���(o��Wx�|���.;a���R4��wK�_#�˙�����L~i��Q�����;��A�-:cZ;+aw��݀Q�:5��DOW�����4.���qb˲_�`H2����搝
#'�;��0�W޴ٷK�c�����+���W����ƭ��u�6��$����;��i�`�^u�����T�5	y�W���+q}N�N�㸁�<�#��*DqT�~ҍiz���=8P+�/�o��odD=���KyQF�l���Zw|τ2Eǒ����ٓ�Ji8MGPNH^�g9�5���7��?��x(^V�N|���S��P��
�S@��'�Tz�M	Uf򘭥��j�2�i&lvT`��&�6;�qu�A�[G�컠#�� ��P�į���H�(oZ���N�f�e'y6�1�Cm8f�����7iɻ'.�A��)�c��0�.��hŘ4h�rHg��N��IǤ,Ň�Yաv�WnxV��O8��T�{���֝�>~s}9O��1-'�%y�E�phda��+K�����1�'�Y�e�C걽�9ɫ��}�b�Ȓ�!�ܕ.r��Ɩ�b�!�V|����I�J��p̡7�����u���=�'/�ł�Ng��z.�7b~i%��b��׉γ��y�0N�尪��t�6�3҉>r��qx�_��݇F�/� eil�)��5����I]�)`G~fL�tld/��N��O����X���^ڑ�s�U��|�|L��Xn�)��-�j��)bnb�(9c���V� 7@ȿ��`v �s�D=���9���,S����	�@�{e�����a˯��2n~�u,,��٢
�wDX�☗;���8FYxt�v��\�g����������{Ր_S3��x
j��L٤&�SU����)�r(������f'_0�2��zG�����'��]YT�@�D�F��KڣfFq�e�j��N����t�9e��6�ˤ|�}HW�<�X���SI�g; ���W2N��c��ޔ�[xj#>�͐�n(5j���>�TҠ�-;��%�k�C�ɛ�W�̿���S饃J7���N��v�S������$�*��Լ���דc15��gǝ��K͛u�F�D�o��R]3�y^4sm�0rD�S��(��IQ:u}���R<N��LBу�� 	����nd�_���C��!'�o�8'='q��.5�+[f"���|��->�u�'��ef[-�!��x�֜ ]����^���t�C�&<���~�D|zx��c;�1��(�t*Z�y�q�T�mQ����I�u_�mF��f�.@5��CE�M�T�ۋ�'����T���N�lmG�����6N�^ĢT����A/�3sq���l��������_��o3G��*yے�D���f�5�ۃs;��j]?rS7�e���ZiB��1q8O]eZ�n�8�\��e�VJϩ?��Dz�.�S��.i;�G��3wh8r;��|����q����ţ�}�Qu���C�9�ggfڮ�����匵�-M�W����d(�L«�����?�$1�M-��Ç�o���XX�� 6�ss��j�	�+�2�
t������i~>KQ�[S�"x]�	�Þ��#|ٰ3������r �2 �e��\�� ��8��~�)w���2M1�4�Fi 8�����aг�� �,H�/�B����� ��@Ǥր"�?d�AM���Q
�:�VI�	��!N����l����t���ڄt~)��։l���42�dlP��m�:��i�J���dܲ7L��`�J�˫�YS>N��)@��ty���S%Yh���a������x��Ob�֝8~�$κ�Xb�_Z��:�������ހmds�5s�	EztP��&ۚ	P��{�7��}$�|qǱ9'���i�m6i�Z~��>�m��8����8�mzSQV��|�it�*�@����in6fZ3����r�N�u���ʻB�ԫ�����.���ؼ|%f���(����x{rV|�#�Q�!�!H;�'��F�J�rlK�H�$m,;�W�^B��筬�K�K9O��֗_��ݻ�4�.������r���c�ܦ���=��x��7��"�����-nЋ�K�� ?mޒ���O��=�<d��&�*Y�)/:׫�J��2���$��LM��{<
�hqTZ�JY��N@S鵜z�oYB[���%��� :�iEK(��@[��U?���-��I����ءrUf�N'��+L�w����ߝ�� �Ɛ�6;;���G�������H˘1�� c�l �C&��A�QApgo�M�ɇ��W�?q�����r������v�<�d9p�~����O�#�A���Rt�9yu	x�kx��8w�1��SzEg����e���NO~h�đ�#���0�9Q����f~Mʓ�A2�˽�#|�A2*�N\���9Q��Q��yKy�|5�d�T#���6ˤ���r�mp��Z�&ӊ'���*}2m2��Ҙ������H>x��m�9+��і|��L�Ƒ.~v��O~��������G����G~>�����/-��Hǁh��(�%Ɂ�_&v�uR��6�@�nŀox/��/��FGpi��ȕ��&b��\qn��H7^5Q�Q�ߔ��S9�1��K
�Q����j�[�[S�Q�K��4?����%����@�lON����76�J��s;��چV�U�IѪ��.n�?�Y���Y�)�Bؐ��<� u\�E�/O�|��n/��<���mt>�����[\���q�w��7䔶�s�Ƿ�F���h�G�Ӎ����;؏�kWbI�1#�m�����9��2
G������pf[�6�2.�4�*��&�����e���'�!��1�J�y���8B�{ELD��I0�l����f���ͪ� �Jc�с3�\^^�c���I(:�g :u^<M����N�_ ڜ���4�����?�CM���tD�ӧ�&N�O��Pӈ
j0���Ȳ3�Ngu�*|ʐ��Mg��$@>t��&@|��W�NH9p(�K�tL�ἡñ�@J��P85E���R���q$qT�;�wB����z*c�[d˶�8�����Ց��H��vTuN
�=P7�8�����)� e��Й�υ�y.ڠ�7%�+-*��P)d���8�f��:P�|N�8���6Pt2�����#�aÓy%�Hn���@��,?�[�
*ƞU���b=��uJ��p�p3�1�ۏǟ}�?�,�oݍ��aL����^�x[O�w�#� ��byu%�ԗ����K�fqĸe���V�*$m̈́��H:��I�F�M=([!/���=ڱ�)n=�}��6�?�U�&-P\�srhu��vc������W�����M�y�2/ ��n?ڭ�X�؈�rFV�]���W��nGg� ^lŬ�Y,�gÎ'�r�b�_�G�#G^����\�Q���H�^	ӏ? �#��2�Ƹ��C�@�5�SR�l��sjϩ^7�<�������i�ȱ�k$'ˋq��ƅގ����C��w�''}��y�������6/�������^U��^�P�%�m@H�T�Ny�[�*,�gڶ�����Fk�Ҧ�&L�xiC5(�yYg�υ���=�[�:b/ s
�[�ʀ=�Ϧa���jӢ�B�#�G: �G�M��4��r�767̟/��I�4����X��w���`�=l�����븩��s�N����WG��i���4(�t���@uh�ѡ0��i�����y�.��I�id�:��'	�Z�ѓ�\2w�٪��E�t��8N�8N��Q��\@@��h��,�G�h�h���t'&>z�n�)�.�2�3p��M�����4�	�̫`z�u�Q�g�A#ۖ�B���;�.�(yrĨ���xM�"�);)
���z�}VG�-�aʺ'eH~2>���V��vQ�������;U`���Ģy&m�L��\@��7�כfu�$�Z�X���|��m�a�Y6�D�V���wTW�/��kk1;� �/�J�<����̩&lh�;62�G��.��8n�t�mӠ�W6g]����nٳ��z�58�7J�iN`99kt�E��`�����W_������ޕ�Վ�ť�[�ׄ:}9i<��Dc�-�em9/��s�]�+�.���r�w㴿�α�/o>�/_����Ӓ,r��*nK[ya`=H�b�������c�S6���2/Ǵl�����C��@��y�e}EG3r��������d[�=9[O�����c��Ř^���һ7Ϟ�����������r��7�[�</O�Y�-�8�<|+�m��Uc3q���M2y%{$^ҡΡ��q�H�vR}���.�Pi�笯���8^8Uf
ڬ����x�¹�~褜<h3y���8��bgx׮]�Q�=Mҭ�:~��7H��;|'46�[ �{{v��L�9]M���Gpfg��8@��f�V��k�<`)���C#-��DW�ew�;�Й�P8'����������Oe�i�|Ѡ<y��eV�E�mh��霓uWg%Lr������&-�8*P�/�qDG��O�PӰƠ�0���z�Ïu�N!��� ��OƢ �%�&��33 ��p�ȇ��
�~�f���;�K���Dk�A�󰯂l�*Kq�8b3�S�։+{��gVnu�-%�I�'O�)�d�&�
 mT�[�F�R��Oz�P���m�䃉wK(y(�c�?� Oe吝��j&�����Z�r�R���z,�~=v�<�b_�(�x��q=��/��ۿ�}<�����!�VӇ��y&����O��FjQ�'?�����e$��$���>�t�i��5t��S�:idy��Τ�qeFN���yl�ۋ��x&���&�?���ї|]Vw'�։���X�V�`O?���ތc9�:V�mčwގ����
�t�����ý8���0ouZ�at?��p���?�o���;����g�K}4L��%�*�s�<�,pKܴ�f,�����յ�+�Ϙ*ۘ�3`�c����X��=��^,-����LgN�lK�S��KKlcy�%<_ߴ�/b/�,w#Osf��m��
�e79�g��q��-]��J�ec��9�y�Ge���:gܮ�5lV�&˺|�K� �س�8���=>�k��t�^�kNnI��.�vV56!i���q��iV�ݖ)�$�I>_�CPy�g��J�_ ����e	�����ۺ�\�@Ѷ�b��X�rJ��R��>i١jK�2N�+N��p ������1�R�5�3
�%'�q>��'�C���&��9Pi�qgL�?�Q��>.�t`�����p]g�^��R�(y �$�r���1�}e���u�x�M,�2���o�H�G�W}�8��'�S��"���m䉜�\�Y�g�t�(V7FZK8��v�Y2M�-�UL����B�-��A�l���@�$��X���Ip6@��t�S���Հi���i���9ꞙ�3>��=7�L9e�
g�bN����(�VD�-Xz��]�nl7�����җӲԞ�Y�s����ѡ���ڹ�17��m	P���(+�XA�~��'x�ll?�n�Ft>m�+�fR��@=3��lo��5��5	
aZm8O�&��G���ǟ��7�F��ǔd�Iֹ��X�8ggeqa)���u������ַqt�K�rP���q7v�?�G�܌ý�vԦq��b��X��m9/~j��*�&8�ǃ�&�Y��t6�߂�P���X&t��Þ_Ȟv2.[��e'Ӏ,�ş\��Nt�����y��{ҏ=��[�7䤟IG!�=������pk+�������b�\:��}'���NcN�/���d7#se���
?P�cʚ�� ߔ��m�iY`�3.u8[��G�~������Έ��~���{����Z�>���x��h1&���������St�ô)m��C�)b9��oS���%͙����G_��@�$p���7������A��ݻ��W_��V$W�ٌ�I'�ӦC:5q��6�B�I�)n Ny���9GǩC�:B�<TG<���c2e2��s����R��SY�"���a�<�c�{��ȟ��a>���G�P����3)+��ק�� WW�|�������<��咔q:g�$����$L��ij���#y#n�T
9�����P%NkYF����ʑ��d2���dw7��^h�=��~��qE�UM>h�����m蒰[��5M]� �����Y�\������2��+pOi��u�IK}��Zr:O%�P�����?'�-s���$���s��Z[��͵�p�Z��曚w{���W�M�������8w�b�-/�\�����S]���=>�3�	��F_�3AId=7�#9u�D��''.�R�Y/��҃��;�?��{���Ν���_Ƣ��9:�'��9싫���3P���"������om3����lo���������B�Nǲ��Prj<h�-ťׯ�����Y���䤞��F���z�]�h?~�V2��ԛ�@�D���P����S��[���ј��omǁ�A[�WZ�����6�>x,�V<��9`�q�~�E�����,^�ko��׉���]P��%��#Ȅj'�cM��r\O^S�����6(S���L+�~��)�4�t�7�Pt_� �2�Ɓ�/�;V�f�-�����jQ���;���:9:�csn�V�s�5�����^\<���xL=�}Y~���xx��w���l����o~�6�y�n�W�v�֘�\�Ѥ1U�g���dXYH�v�8w8�vT���1(�11�IpnSftU�8a�Nw��Ƹ?����y3@�n�;E�8�:�r\�5���^����	L��c3�-��b^	���?��&���'h{��e@_�]�G���̫:qX����
N���C?u�Xi�0�\�����48�1*^up;[��Q��!� Ϸ�X���;��n<��xz�ft�>���0��r�T���Hε�-�<�L-�`� sOJ��s�"����N��A�t��m"\��*T��'�h��*�	+.��[x��^,+�}ԉ�_}���������X^�������2t8OlEp^���nĥk����">��x�h:Y^�P�����^��c��VzAܮ��8�^�,�_#�(�l�:������7�R�e9�٧�M���M|�Obn7V������ν;�}�(�r�8�m�$�����b^c����x��ױ{�v��ykɡ�=��ܿ��0��<���#9$=9Zm����R�_؈7�����q�_g{Gq������rd',y�����U�>r�1 <'�L����IYI�sp��ҹmö-V��t��=:؏�t�7"g�h-HŇ/������ُ����х	e����W�]����cjuUm��ۣ<HV���!��Nr|��\�*�Jϋ� �F�P�@�V��\�~�:X����������u�8u'�c�@."�sn�u��%��c(��b��V��\Nxv�<6�:��x��d_��F�C�;���SZ���N�_���~���z�����ev��[7��nE���Á��Y��+5xega�S���e�K��iS���u���hAh%�qG�4n����)����GlS�ҫ.�
��*�V�7	��%8���,P�,� �ZvG���i�"=��@��̼���\�����jK�h_�чy���Y�2NH�n�.��VH��-	4�`�����=���7oǋ/�����1�ڊދ��[wFgw�u�x@{��m-�#қ��.5Y���
�w�i�G�n��TP2 %7 Ϻi�<P�����kϪN9a�b�27-ҝ{��G�ĳ/����m9�3q�ʅ�b�G��4A0���窆h�ε�dr[�wwv�x�	f~��;��J�꥘]Yt���x�}F�jnca���=�IHyR��	|n%���q};Rc��
�%�I�@����}N���9���wc���=>��t�Х�x��?���n��r���d�ā��x�4�xS��(��x��;�3���X�,���,'�g
w��sON�Vw�Lozs5���4W&�ư�|��9�'q���~�l�g���	.������;�&��J�%ۙ�3�(���q(gSɬ⭨�y��[�=]�,�����@v��gS��Q[l��f,\��ggٴU��r��'��PP2��d<O�;�I�82��-H=�xT~�$)X?
.�M><XU�d��~�,�.h���<�-��>'��Q0?�q�l�U�Օ�XYZ��c�I���������}��;a��^ħ�~�[�\9b-E[�%�R���� ��{�b�e��'�\��( ��f�k����f��]��i��W�� d]���7��'_�LK����y�Ьs�85y�ySf*�qg�3����û�y(���|�=�Z��'�׏x���L�	���y2qI�CC�r�Q���H9��q���_q��7}t�_�;o�=S�ŀ#H`��3&p9N��Xa�g{'v��6BW��;��?8�u�ǖ���8�W�tcfq!V6���ڪ��ȺE������?^�������  �	@�^��%/`�H�2�[���>#�g85��4Zr8�?��|�>�"f%�$�;���l�^��PK�p��^�؊{����e��AU�:r��^��ɯ49�|�h��F,�ߌ���&[��	[]��r<���՜���(Y�/�*�JK��g8۴3�#RL8�)���Ⳇ��(}�-��N���8|�X���G�1�c&R3����oąދ��fT�%gj��Ǐc��X;�z3S��¹��9M��W<�?��������b�+'rF���"��4��7�R��~�#e��9����IG+ǭr�o
OX�O��q����RE�fP�.X;[�e,D��0��0��������Ҽ.���ԗ��ݕ}PL�1o���46�z+��^�� �����l�q������xr[�p\tF�.\���C���R��7�%m���~%NF����s��+/�stO�m�<.��)M�Z�7#ټ���i�f��L׿�ۤ�9���ݤ|y2k�k�t�i�'�Ν/(�����2��w'�`��<���o���g���s�)��Q`r	}[���fWs�3)�UG�\�`�M>G.���;���v�5�x S�:G@��#�+Y:�As�-��X_)�g�\�|�ï:Ǌ���>PG���M�ˈ���H�@��$+=����A?Θlu��$]�zc�%V��'�S�Ǻ}�=18�`�J���^q��dFʢ|]���y�d�G��'d�� �\�l��@�*=YǙ��0	ļ�bM޽��J�X�W�@�fcN��8�\������X�X5zO��~�Bס�^?��6��c]�z�#�����X�X��y�<�Λ�����џ�϶	3*f��L����lQ���V�&�jc�<�9�z՟'�{��>1�� z�Q��wb뫯���~���Ek�7߼U���bva�Y"��ܽ�>�cl�U��ǹ�v������gq�	�L:�uc��iN%s{^N��X����Ԣ�Bu�"J3N�����8y-i�,^��!&�W	K��ɟɤ�D�}Nz��z�S���7��>�!O�ؑTP|�Z��S�bi�'��Cwg+�?�C9���0�j��\+�/H�����^a���>{��{v��s�|�y,�}�$���ݑ+�}�to��ã���ۍc�%z뛱z���Z����Ms��L��͂Y�;��+WR�be�� g:,�&��@���/��N�=��o�r[�-zaNN��j̮��i��]����|���Dyױ(�����Ôt�&�j?�?��[�����H�vkA�T��<�4T��xa�ϕڜtڍt6��3Cc"�dd�H�h�ғN: |r�D&��1����$0�O �ǈcK�H֭�a=�Y\^n������]� r�=��m ��V���b#��Qe	��i���B�E�38pn݉h���"��.8|l�S1/C���� �����ߝ0A548������_���g�@>� ��cLf�1t褡���⾽��xQN?p�:��-�1�2�2�2:߆hdc+;W�������xBp�����
�C�r�9N[�;�ޤ^��Y#O3��0�ϰ5#ω���N�ϭ<�����Ǐ�ٗ_�ɋ�����El��d�Y U��v)7�+ �j�>�
��J���p����AmA����#H�?|��p�g9���xsD
��mE��Z3�k�
�~��N�9�Br4gxCx}�l�_�@�&�L6�Îmq���8���\��������h����:��d�������W�:²x���l�MB:�>F���8�����)��+Ѓh�ԏ��l�v��a=y"���o �_�/���ƹ�W�$�ĳ�7��_�ӏ?��v�����{�$�Ϸ}[m���wscV��y]@m\�/]�����-UyC�Ejr��������yQ�lvaQJ?L����$�}@G$/��]P�I#�PS�zɴS��8�m�ʌ줿��O���	Et���� �x��)[��F����`O���pT`%�la.����Wg���W�T���fVcSۓ��΅�ډƫ��F,��(;�K�^��[S8b���Ɔ�u�r"�d��/���@�BⓆ=U:�v������q���#���.��mƅ+We��_z��d�7�Յ�B{���t[��X~�z���f�d���'�GӈwIG!�\���d;�G�⌁ϊ���n��?�
q�T�i#����0��
�GY.l��S�?.�U�N�t�Iv���0N3��/�˶u�9-i����4D�q�ǃF$ �Q�͍��E��ǩ��� 2?�o�w'lX�
(���>�'�V�V���1y �Wd�Ȕ���ǆ�|���1�V�:�&<�F�'H:I�|:Pi�)I(�4�T�
�WPx���bN���㾌[���
� ��">A���x�OW�Ǐ��ǟų?|�������O_������޷7��Cƪ���'j��<�d�v�'��'�*��V�:2>ψ�͉�A?˫��%������
��.uD#Lt��+o��$�������E�J��??=�����,��.ϯx5�sx�/����-�kR\��#9 LL *t^�t)�WT�n��]��l�؆�u�O�du��NQ�$����GP�(��Q���%}QW �p
Ix8�����{�(zO_���'v���x�4�.]��׮�څ*s��_���{�y�4ZG�8�?���nt�n���g1�ڏӣ#���+̷c��9�!9�c����x��\�]Y���E߮9[�R�W�,�x�6؅�}���G��-���*�u4���ūG6���`g��H����n���Q��#��%�=8�]��e]����V<�s�U�aCW�t�߅�W������JʱK��AΉ�!ʆؓmvf.��m��#^p��xSU?���c�L2NiLc[�r����������c��Ԫ���C�e{I}��6��Q��EsN�����1-��D�CW6�].Z|!�qbqF��.�o������DOeg�f����mNː�	!��",�m� y�c�閣)�l8��V�W˔=!5�E�&���g}�R���Z����[��Xu�I��]�}��k᧾ɇ?�7�HO{f�缡I]J�❕@�SW@�R����]�!��k~���l#�wB�3Is�����	L64�������o~�뱨	φ����v����1�W�h�Af�ư�vz6��&��c�е@����F��50j���$x���W���.¨�2��+���Q�d�d|�(n�C�|㒦r��j�A����:qt�Onw~��ؿs'ښX�{Gq���=������k��D1�����rR�WWR�Jg"���f�c�*� ��� l�G<�r"K��@&�(N���>I;qFGA����M�8���I�Y]�N�ĳ۷�܎Y&�����2�I�D+t:��<w�W��/�9�665a�DW���R��&%M(r�f�}�����v�I�N����״/&����@L�M�����
��C�j{Ӥ��2�%�3�5�d���ח�8�=��+�$�+��z�R��ӟ��;o��ƚ����?7�{�'/bQ,�HG�?�m�����]����C�̵�Nb���غu/=��#��bqmI���ۅ���۔tb����C���#m�<�1a�~`�,��l����F���IH�P�pYUAo�`�C�9�m��N�bQ�?�]�y}|�n����8~�P�^�����n�]�t���{���W����ُ���#�-���L�ș�?6ѝ�?k���l�⹸ �[�g�$��cBe2f�`�Wi'���ps\�8G���F�:˱&�1
|t�:J�6'p1�8�)S�ԅS��N�Z�����q��[���/��4|��a���@�n�N/�ǅ�|�E���V���\ ��J}�]�KYlCF���O�/r�.<�drO�㠿�x�%�z���C�	@���1]��y	�W �?�lѷY��À�.�:�:Y���>ن0�<�펌�KYn�e]��Eߋ	�_Ը�#��{��҄��3i��/��&(c!`|��8::������Cپ�ؔ�n�pr�q�Hz��hl<U�A�V���X'#/�7`�#�t�"��L�ʧ㛆�'Y�6���P&�(� �@�Qʢ�F|*��	%�� �Ab�&]��ĉ�S_��1�P`؏~�(N=O�S�A�g���d������PY�HG�_z����<<��&�Q{���(=Q&��
�(=Y�G����S]q���(�ǝ�?�����sq�����Ң&��Jg�<1�-��}+|ie9�_�
l8��U{go?���(]����܃/]4,hBZX^��ZOT8��v*l���3N���5���(>a����[e�
��Ky�'�Ձz|h��F�3��vl!p��y�nŀmz9���^[�Ko�KW/���Jt��r����僭�<ێpM'Wx�x�
{���·'�8���aL�qa#O��R��_Y�ٵu�t��+>���~�!;�Qr)?�Q0���<���/�Ƹ脐iP�Q��WPZ��od�"���ON�D���d�K '�1}t$]��T��&m����߂V�?x{��ގ����^�`l��<�9��!],��T��(�]���_��+���ؘi�b���q-^ie;M��x)�1}ב�}ۑhl,�#�T��Ѻ�.ْ��i�)]u�M�4�hL�� ����ٽ�����8|�H(�r�z�P�m��F��� ��X{�m���&�S]����Gm�|��kB�蜴�14W����ej,$rI&�^�Ȭz(Cv�q�p��C�SG�&ngPe��-*O�
�8wH�\� s��r��c�#��r�'��:�����иp��Ɓ�i�1�Se�����	hW����v㫯����"��{ H#C���~���~��~T�����FI=:zrT9�a��+c$md�ԱB�[Ց?�� �!�NIC��te��&p�Wj����}�z=�x_��ܰC����M9V]?d~��P���`��d��þI�R�L��o�!�PyVR@Cgy�M�������fb������ Z� ��5EO<�ul��6���b��v�J�d�>y�_�>�"N���X����R,����#屹�N7:ҁ�Zh�)o�]܌�iMܞ���w�؀����B̟یs�݈�Ғ70��)�9-n����P󚘘��q?C��{�3H$*�8��t�^�IΆmS	#L�B�~~���y��4��n������n>zbg���g�bV�N-/z���tlH�#���w�#��_N��7ϛ��K��}�<��IǬ@����v8���r�:rNfV7buy�����Jm��ccGt�b�E-��M�Q#�G��~�8ݿ�P��9
*~|{F8�5���w9�ǻ;1����0��9��tɋ�<K�}zO=�#�'r�pDٺ�gQ]�~vV�/�����.l:�|��o��ո�_�y��pkU��יe�>��ѓ.�b>tM��Q��r����@���O@?���5i��-(�����T+�p����/(�A�ї��7���qz�'�
��C��o���Ӂlh��7bEaf}ݫ`<?�sry�QcG�H��N�Qr���@^�}e�S�h�(b}�W{���Ɛ4�v2�qt��Dۈa���87߮GY��2.�}���k���s]�q
�V��,�]���A�۱׮]oT� ��3�W�U�$������� hV5�g�}Ϟ=mV���p#y,��U'�W+c��>�u:iV���!nCͷ�DJ�NLՏ��9�28�ԏ3��c�����DG�B�_����q���vh��mg�9/�E��9�z_�Y��ms%��,�[��s��L��X�8�	�ψ����8����V׷��[ng�~L��%^�چ&�%�3�:W��f�0�Ν�Q��3L*w�������T��v�� �聉M2M�L4�t���ԉ]E;RÝ�ؽ}/���۷�D_*O��j�y]�Ϯ,�5�;�S��/���}�ciyA=v*n�-���At�=�]M�*ϭ49,���X�r)f����wc�%���}@Y�&$����B�Z�>��X^e���Vu��8� ���Q6a=q�9W�$[7;b䫮!��A'<,~p]ɲ��I�4�*��@_�[�9�-�<~�<�U<��+9����gy�ŏ�@^;�3�����*��b�߭�[h�6��>�6�ϝ����8<<V�{Rj�b���D'�6]�A���Ș���A:,�#�pSO��+��vprpz�E���E��}ُl��MoJ��[�1��An��I��jwn�!����A�yɂ3Ã�<wy4?3�/ǵ�U���O�(@_vϋ1ܮ����C[{5Z�[�r�7 '섒�	�N���A'�?���6ob�t�9[��gۈ	���,�Ѕ�l�LrS�������ؘm�š�����˛������[1w�b��ͩ_i�쳺ȡʲׂ:�t
��}{���J�9�9!�
eh�t*ٝ�<���Pi�%n#�`\>���hlcJ��?�IOno�����7�Ӓ[�l]��8A�A7�lc�Oŧd�g�H�| v��m��(O`^)c�2��Q����u��;%���/��=�e(����N���#`�����4�j�[ZLCP�1�1R0����}�؆�D6��j 	��F�4�b���s�<����
Hw��4Ʀ��FuĬ����=A�A8�g:M=�4q��k:NI ��
��*���&o�͉ ̓�����bn^W�H4X�m^�W����j���UN���%�:���+��<x��d�����B���)SXb K%���|���H>'���נ���x�	��N�%?�ʃm\ j;�hl���G1�l;N������ѕ#�Z\���1���f��vt�||�m�~�Ml=|����V<��ko�0ųa��$���Z,nl��9]�5����ّ�6 N>msVM����0��4��*�j_��wJ�FcϖᝎNHO|�����S�w���IVzK�ԡd9������ễG�{q����<�������u�V�n�b��q�j�]�EӍ7^�������±�9M�t��|yCΊ���)�n�Gg����S�ަ�zx�5o1�l
�M3�e$-m�dC��7����9��7u�3��^@��%Ӗ�Y��
n�����0llnĊ��@m�u�o�٫w*N[ٱ��%yOp�6���달h�>/ �!��q�{��/�����Kq�>�7���1snSz�D>��������vM��}��\$[TAÆ��(�_��"RL�0P�����G��q;�||:SjM�;� ���{]t𩢣�8:�đ��[jŒ�7�x��?��1']N��-;�I.���KO5���To:_9�慴�~��E�B'�7��*�<'�2��a�uޠg]I#�I(H�5�z�
����ҡ�q�(K�`~�֐t����Ǥ�I�:sRޜ�Lm���%��F@�o��"ں��f_x������T����0�q>z7o~+|��P�38`�6�ƠI���DZNn$���[��k =����FJxŸ&;��9�	� A(�@�'c�Icv��]��q&�����Wy'�j�P�w<�C��1�I�}��_���~'��40�I9z�"�݁w����r.f7��L)�Z�� 6N��c"1?fC��+��M�_f��c��?QVG�҉EΘ������.�399aS�qx[�շwb��C;U�p��
yf}%��WcF����Bl��8������O�-G�Ӎg���ѝ����oKɫ�
���K�+�h8�ߍ����}~}a�6#�?���6�xͻ���f����
^j[������%4qN؞�@��{^T �G`��Ԕ=�P���l�1��:�Ά����gx�r����L�r�X�c����X��G��ۛ|���x�m�O����c{2#��mM
m>0,;�/8(B�Lt��䄹]�8Y�����w���dgV�5Z���F��_�S��P_S�װ�.�.�����l ���h�[�<�U������S'��-�d�.�î/~p3��''��c����������X|�Z�v�g�WK�	�y��{�M��o�I�F~�EL�Rrb貜.Fv"�	֡�3S�X�=0��y��	���i����r������a<V?X|�r����x���[��~���v��X��C�L�Ǒsl^Q�E�OB>���Gϲ5V��qI�O���A�o���@�!�.H+',/�g��-�(�ͱ�{|�q^�#<2T�΀ݏe�.0�V)��U�C>����y�]`�L���l���>3�2 u����	���0L�:�������S9a+^��s2��|ʌ�|������`ԩ��K�y��\��)Ϲ�k�� �W��x &@ٿ�U]y>��T�q�xA:	�f�%n�-|��\��<�L��K�AX'N{����i��X�#NYK�♖%M<�ӝD��R�̶�=<���N�i�铘]^���99l��4q+U�P#���=XpTq��(�|*����\���.���y�9!����loH��
y=�*�ae���&���N��	������l�	c!�/_���_��k7ba�7=�;���7���QLs˱׍����l�����N��)���9�6�����{�u�V<{ˋk���	�'[g�g� .ޙ���ߚ�2ql�PJ'�'�㐺An�ʹЙ�EGj{:�`���r����cIN�p�L�ї#v�;�v��@s�׉��}9�}�kE�LK�Ў���p��Տ�C�&p��0����Y�G�=Ւo'�4������+���+�/���	�#퉬r �=�u-/r#g���@�ϤӲ{VK�:�(W4�M�4�ϰ\�ck` Z|+��[oǍwߋ�t�r��5����=���Ab�	���h�N�py�g�L�X��{�'q�n���q�g?�w儵���uy��(V�ǜ�¶h�b����n'O|��]D��q2̪�Aˬ�ǺI�(;�@�V���*Ϗ(������c�U�/�4o9�l�������H�����G���'������Wq狛����x#��#;�N"���r(�տYU|y�˘P6�m��&)(蠃�|���4���\Pz+��Q�V8u灲�3�\]]����8�������|W�W�-���l�����(y ��H���.^����
�V�
9����朰2�#z��~|��cY�WS {�0��&"�#�Y�$J��$�c������g~Ӂ�NUFm>��Io�:׉�>�4�����I�@�`����A����Ȣ:+��}l��_rP�\�`��AsFW�'/����B��|��[1h����������I�;;�ś�g�����<sD�����&C��<Q7ϪT��|<�b��#��x���%Ph@�"�n�[ϴ���y�7G��q��G����h2���^����sq�����[����F���hHO���}���xf�bZ�)o��t�ˤ��$/�73s�8ӊ����g����S��05��kk~�/\V̬5
��X^��.$3��u�$;!��r1 ���_�e}46���Թ�'z���	uV�D�z�3�tnUN�<3����=��������د�h�[��p�y�ݎ��|�Ȟ��+"8�r��])O��A1Y�lv*�dQ��6�͟�"��\���-n6%�eK�ԛ�*��41��M���!Z:_��2����H�,Wz���
�~E��V*�NTG�o-.�9�ͩd~t�~l?z�Bo=���?Y%{�$�`���������ac���B+ο�N���_���C�a�ҵ����ݽ8��(n�y<�wOU�u~.��'��_�g<;)JO����j��e��t�R�z�q�&yt�Ð����GA(����L���O�c �<�6/��ۏW�{#�����W�������퇺 ���~��JW�ؤY̌ [��g�+ n_:�"y��lg��{��@_�?QU����d�p�,�Я��@��-%M���i֝�N{;v���{~��3Q���y����EdC�ㆀ�����UK�s�&o�����F�������A�C������#�90䲜��'���mV��a�P��q1��A� ��ڐ���W�B��Ί)`���v�uũc3���� H���SƆm���'>ىˀ�"�|	���XuO��74�V�<Bu���ͳ��v���~]o�w����;oƝ?�N�� V75q��$^ܺ���u4�ȡ���R�^��.k���S�7DUȓ�&��3pV��mIc��k�U#����<���{�d#]�v:�K�C���I�2����PNX�������Mv�����X�x%��c�x�����غ{;�:G���g�=�T¹�W��99K3�8=:����{������8�u���C�srreӼy�^k^�E!�����[nJ��=��x�o�M�M N�(oM�Sp�&qOl<�/�Q�iҟ�#�Ӓ>Vc�%'�t*:J?>���I����C�����N۳r����v�O�ZD_?�C�R�'S�Y�u�jGG��ե�������~˗.E�5�z�^O���?�!N*�_�%��D�3-��R/�f{`L@g�'n�V&Xq#_?[��K�)�'XՂ����8��������G�'w��L��-*p��Duv>7_=�낦5��|+.\�1j�����R�C9���y#^��r�ݷ�G�Ԕt�zv�݌޳����~���I<��Vl=z�α��\,o�E{i!�G�Ԍ�o���od�+�[���@��x��L�s�HG��Ц]HS�^M���	k�ƹ6�I�����]\�S������{�,�s+���GO��-�����Qk*�bgF}�^��8��<0�|X�+ػW��x��vs��N7�͸�#+�֏�!��0]3�q�=u���?����:k��)�/�$?5��\��-d� �P�;�C���:�7�>4M�F &@�Y�e�0�S!Ә,�*$O97*�}��9'���TW���s����o��`w����ꐱ��'m�(��-+�4L�.�u��4�X��G����/?�ҘHH��O˝*tL��,���[H�|��L��W���#2�W�[���2xB��+>ɏN��u _瀷��㪜��5)�=�Hm?�����|���ęʹ���I�z���Q,tz��+��~G�b,i�?�|\��sS'1�y����+�ظTߓdՂ�l*����h�p��S:�yR�Dq	E���GG�4�+�Ӛ�fO�������e��5<���Nty�Q�ʹ��4i.���s�~~]�$�a7N�o���N^Ġ�Yr����R�����/�9j�T��� �t���F�������m,�&��ʆ&��)O�t�t���hHp;�#=5�,�d'���1_)7�24G�|�.��*óI��З��6�T�
f���^���sq��*'k)g�q"��k��[�3�k��[��Tڼ�,���V#�	���~fb�l.΄w(o����?�k�J:S�_��-Kv�?�� �������G�U�72kO2D�ʜm)������?��DTy@9��}�p�ʹp��S!J.�?��)�z�C�{��(:����C��i.+Ssq,�d�7����$�x�Fܿ� v^��b{^�?�N��A�����+�bcM:?:�[��o�����;���8�w?�Tf��t��֑��F{m%Z�p�֩�!tb��������	y����˾�>�����GӐ�x�/{�^j.���fx�@<II-�ц�Aϫ�3����V<���1x������?x/V�^�����o�K�R�p�v���ƬB�2G�N:F�sE�x� ��m�
��TH��2"r1PZ���_�+e3�H'���&8�=��!������u�{�Qiy��jױ�c���}�b��|����oeB����s
2ӗh_�\�O��������;}�q���΋�I���v��|0_���!MŽ{������B?O�]��H�R���At'�i�i��(��n���_���VF�=�W�ҩM�
�ى�)�*�7���$��d9`��*L�֠@����q^�p&i3�����r�/��w�Fkw?Z�r;x��4�����������0w�� ���8��q�ݺ7?���;1��+���o/x���aUw�A��>25-��ҡ�s:�U��d�p(�s�<-=x�%%���D9'��+�U]���i���ȩXo�Q�H�le�,9{�;���ޖ��[��:�`tfa6��&e���8��^&m��w]9�]M,lT1��k�~��B�%ۍy9�(Sۿ�2?e����Z!�L� Y�~���6p��[Z��M�	eN���r\X�k˫v�˔����z}�j��ţ�%�Y`��@a����DT��v;�����������~�O"Ͷ��-�({lɻ�{�|�h���m.T���^ݒ<M���
�?����P�^E��ic��4ǝ�.9���������f�,i�����{/�]�@eNվӲ�+�?�����،G_/>��LXO����rа��Ƴ[w��G�ŝ�m�s+:��rb�d�޹�.^��[��k��e������+|�F���_K�)~ʎN��N�S8؈�'�N*��ǝ�w�)o�"�|�K��{?�|�mlݹ�{��q�2o��ׯ��Ҳ/�k��"��n�i�0�O�T{�G߫��h�N�Q�S�� �	i7�G�t/[#�I���д�DZS��N�R��72�O�2�t:�1A���M:'c�&�t3x<Q`1aMc������2����>VF�Fɪէ�~�I�g��y�0;b6��*�0�Fqҝќ;L�(m"T:@y:�E|2��1;�,M���D��fO��k�+ 濡�	��t�B�S����%ڜ��	]�����q�)9�pM Jݗ�%�k��wxtGݎ����P����rx�Ipg/��};��PW�ᰧT��
&O&l�Q���Hx�G�p\���洎�+�Lc��L̊C��x�ܪ�7��Xaґ&gyқ|�]�c�-oyLё�G�b�֣\�ݭ����8���֭8|�(��<��Q��iK����j���[~F�'��y!�58�s"g�+s��/}]�Ʊp���8ր9�*�F� �������,s���]9�-�a�zЋ�a�ħm���vg�_��A��j�d�х��Xk�Ǖs�cYNԼ�u���fxȞ�=�5+^�E�)'���6��4	������CV�/l��{oƹ��8O�͉X�mL��1;�G_�Ȧ�;w��%�9������ɌD�&d�,ȡP��h�b�Xvt�_��r7z�IM D�&���qh��X_Y�ۏ{�p�����˅������ŏ��Xh�Ń/���_��f���dl��C�r~3����Gq����>��o���a�#⪅�xi��̆�߈����ɮ���3�l�<����U9�@Ʌ�i/)C:)?f�L3(j\����3�с������W���؏p��_
��~����,tdW~�Al��Z�y[hSi�(�[�n�m�
��}#3��?���C2���j_B��<4P85��K�ٰO�I:ƛH�tƴ���l�L#�q�<�&�� ��M\��,��f^��ưu����]��0�����ݎ����EG��ފ�?�<�e&< ʲ4C'vDe�ѿ�靇e5xH+æ�L7�_���Ց� ��<H)I4��?�vi����@S�L�С�i�ī&�t�dZ�����r$�΍���`�!~+(�*��~��
>vv#4�u��!��"e�A�_<�#E����w�?x���G�:�G�+sձ��kr0�����p{BR4��3��٢ ��/������D��e�!����=I(�uonM��j)yFG�c��[�{[ےa'Nv�bNW�xve����S���ưs$�|t9����y�6<֕�:rX;r�p�l��\�y�M0]�}*�f���ؼz%��V�ê]~��rPF�;i��dmÚ�\@P��4��.�6�<���Ʊ�s��;Y�c�~a��ߋ��O�pK:��y�T �)g����+>�]��/�~��q*��r�6�z=6�|=6_���1�7I������G�b뫛��/���bue�on�L�9�f��o��"�/�PM���.�vR2���TA�?�������2@�繬��_�#Ʋ��t+����.-�k�,���'�$��7���G�Fww;���Ԋ���K�PV���m�p{/N_���q?V$'����:�ln�tU���ڬ}*��l&��]�,�Q�����`��W��trG0���eZ-;�#g(U �NN��M9ry�u��\r��x�~){ns�o��)H��o���ok�nS�qOУ^����Wg�O<Ќ�����F�;�뎊!I���N�)�sꩺ�����U�:�SY;AM9�iHS�I�5�/d�d�C�#�,t��ב2�[�YW�:����С��$� �2|���Q�X�X��5I��%��{+ajtO<jC�/��"��I=PƃS�j�O�(]��t���Dp��f�	�N��3!�W� ;d۸uh��obd�O9_Y_�R�<q2�H/^��x:����yC�W�����9�J�d�A}�����N�>��� �:���p�u��n��
V�@��xQ·�ԑْ`A��<��4a�cIN����WzN[�59 /�a��C�ΰt��'X70��]ñ|ƶ.ѡ�3+�sdfP�l�4<��'���i�Xb�'>�r"r��NL���C�!���r��L�Μɑdb`�\�_>���D���E������8-����_��"'��*{c3��������j��L��ⴰ���%/Ǥ��m\�zh��)}MB�7'pa��ږ@hppL|�Xi�����[q����pW��0*6�օ��B̬,���F��~5.\�3J��og���T����y�J\�r-.��m9-����c��8�ӻs�n�޻C�8��P@��k˱r.ou���U߆y�k��-��}p�$P e�N�G�����"�1��_:�c��x�o~aIc�It4~-�ĵ������k����x����}�Զ4�7#¼(2���� G�#G��B��s��zy��[�$O�Ȫ��$q$���B,H�׮��
�+�Ƭ�1�iE
X:������W �یg9���}V>��o��!+��$���H�\<��}'ο���5?o�ŷym�.��P�?G�CE�򠖔{.B�:�`�?���/ھ0ױ�)���jH�#��]�ij_t��sU�s;��3���*[��~�]�''e�7OH#؉m��B.�!�Y7oH�qk������D��7�LX}����~�or���	�0y�φ�r��� ���������p�,�����j�;(�Y�c�G�(�A)��cG�Μ�&�&�v�m��iz��&;( M��䱠�MO`�$3u��U�ʁo�G糬 �C�&��8a�'O�Y���[1+�+o�Ƿy���r��VW�8�G��gU�+=9/�K��?:���g�WcZm��U�k�3��g���9T@��tl�.�C�˶|��G����\�^���p<o��$�)��)h]Xٌ��%{>;ۏ%�@�%�\/��eB��!Ǭ=�v[�o:u�]��I̲�OeU�����EW���;o��?�y���F�.����G�����Ń��6"�o�����}���϶n�y�I�����a7�N�s��n��3h��N=�+~${u}-XU���R-*ߚ�c;���X�zYؕ���uZN���n���H��nQ^ք{�굸z�ZLu������}��/����gxqb�ۉ�5�1�ǋj�9���ʚ���Ǔ�xd���˃~�&r9'�X����7'��u���yҁFo��v:=9�n�.�F�]�o��j�Vl?|�>�"�}������.̴䈩����^϶��ZR���,R_\2."fK���S�Q��;_]���?����ױz�rte.o�Mq��e�c�	yR�S�J��$R�Y�2�@Hg�t8�=�ې���J��?�hټt!V/��˯��0�n����Z�	��	��<�Mz��Y�j�7�ߔ/܂*Cz��,@���s@��y�������~��	�f��x�y��.����86ȍ���R�؎���?s)/.ԭɜ��#t0�\ ϫ�k�I�q�:��d{�.���o�	S���,���������1V��l�1�	HMC�U��#K�ixi�#\:�N����z�ä�D9�6��J�Gg0:��ۑh�W���
8?w܆�oa�R>��S��%��4P�E����#W5xu�DNG�h?���ܽ���]n?��kY=�o���a�51�b9�У.V4q����!~���ך�}�j�ܹ�Y\H�O�NN��-�r�)����br9nKDB����z*]0~*!��ѧ
�� |�
�S+܊�! g��꣥�R�I�a����vt�M1Xf{�\��ͣ)�C�UYt[�|҆7ӈ�e�x4�yJ�a�}�5�C1��kq�'?��7^��ԕ?Ω&xA.�|Pq�é� �x`����"(,Ӳ8�3���LN*-�x���Q�E�`�j"�r[G��`�o{w/:j����wߎ��\�q=�������HNn;n^��U0��T����������;�ݹ6��6��+[��E�#��QG�b����%	Ot�nO�b�B�p�V�z�s� z�gg�KuaD)��ˋ(�-�E��|#��К��~�h��>Б���WT���&}������Oc��0Nt�3�Kl#!�v_P����ڶ�h���M��ט��V�����;�����rd������O�z�j��ƾ�d���y��B�l�t>	/CcG���3��p ��K*�>�x, ����|�hVA�Lp&G�D��?��AurU��UcG�F�>��)��?��x:#�8������
c�gP�'��Aؕ;�+P8ֱ��(h^�$�9�T�肿��M���LQ�s�r>�:�"�Dהx���<il}7cG��c� �<kGM�����~�&�����s��ٱ[�OW����N��(�nkPR�ʎIi���� 0����cί��p Ic'>P�n��1�tx���Q%Ek\�$�k�g9��2�Rj���?E� �l��:t��$R.�O�G����������ǩ%�Tvw��ރ8y��+[�Z-�.����`��� 6��\Z�@_�{� ����@��YZ��+�cI�4"��Ḹn�H�A�����'j��[�y%'�cg,�΄����#�� �zl�7�fu5�bw�e9�|(Y�L
�9�\P9M~\��PϣO��(�Y�LԼ-	�����99o�ߌ�� .��N�]���)�hТ�����oo")�����mc �5�G�V�����@�H7.�JG�0ţ_�snp��v~(��K&�y9D�nfuj{o?�kkq��7���ߏW.�nz��A<}��Nk[r�yc�_WX�_[α.�Z^_��-J�7�V�gW�z�1x9��X�<��6'k����������1��C"G5��j�
�H���v	#Z����&_�G��^kC�?[s�={;�ގ�o������6�i���EJ���H�u8����,�r%�/]�͋줰m�ߪ��8��3�F�&V�ׯō��?ǻ����Kd�S���T@[�l�	�5yFF�N�p}�30S?�|���� ���M��ęP��'h$���K7ק ]#ϋ��x�b[|/�������1��n�q�q>�0��u^��AZ�)N���v8�����>��.r���r檎�)y�a�W�,4(;l�w�A;i�G.< V׽���uh��u�oIS�׏�j#���Pݿ��ԇ2(�6u����sP�-9���o��|�����0���k�
�ʀ0�2vw䦣L`(�j������~N�+���W��'��#Ǐ��)�����2���q����Hid�[rY�e��Gz�|�#w�Wp ��6 �>
����L�'r�N݈��8�s/O�ǂx�&��q'��?����|���
��Ȫ��B#��8a���������x�͘b3WM:8a�J!%W�̗>W�_B��L$U><)�!�P��I������R����-VZO�A��ƕsq��X�x56�|^�r5�d�ǲ�^��o�f��Ӛ�D��� /�{ia�G<i@�a�آ���bCNع�_�9%8�􋮈�4��tu>#^�Ս���`6�r���D0j���Ʃ֕!�H������W/r8A_D��&�t.$��l?Z�����cC���r%��xMt#���Mܻ}+V�Vy��9��E�%;���6���K����_�K7�ƕ���X`��0�[C�9S�q[�71y�h(�����n�0x�3~f>�H�-p$��:���$�9�mL��)Tg8z��8Tc}�~����m7:˪ڐO[�޾;��Ǟ�=�O�Q�j`v�_�z1�~�N�x��X���J����98t��n���d����ka)�^{-^���w���K�ݸ=n�N�é�l�7 ��:,����2��4��R6��s�l�W�ʐ�Ǧ^2�(��[��%�������'^�^^�۪���!C��4GE�Y�[�ɨq��zK��p�\F�?��3m�*FU7�=GT�tS�B�0���P�)n<䚼��~��&s	e��h�ʕȴw�T��i�U�a�o�'��_0�qޟ�'�M;�>����H��ɓ�q�ΝX^Z�[J����`V�W�_�Ɣi*㫇fٚɀ��Y�G�$�7�Uw0�h���ӹ�T�96U�65�j ������$-�u^W:�$�5u���C��I����]���6)��T �ƷLTϞL���:��b0�κ�05ɱ�hoJ� �@��e���[^0�>�f�ҷ�T�@���M*?�Q��ᇱ�����X�7��I��d�*�0,cʙ�)v��	�A'Y��*4ns�� > ��(�[$Ѧ���Is������Ÿp�F\�|%�4ɟ��Q�y��/�xsL>^����*��|KN�\��?��+n�Ao=V1D�H���kq��7��59�=�%� � ~Nw��	gO�������o��(��D��'!�F��#�� �Qi:�����ʠ<�D�{u����.�>�N�$kQ�I7����{�����v,�a�p�j�nl���~���K�9y�����j����.��t����.�Ջ�ʕKq�ڕhKk뱴�W.]��ciV����j�g��⶝�ꋯ>+Ls�h�R$'�9��чR/jO��#Dcl������	�I�j��b����Œ���k�)�6;����Dr�){A�-�ߓa?:�#�{G�i�w���b�ꅸ��w�'������~*ُ�ѽ�����)W{�~�Y�{*;�K������?���p!������mb�\=-N���O�/�8·6a���x��tI�xt���J�I�s���B�v�|�M�bO=����X���s���<���{�7i�Ie��?Sw>P�R�e��ZՇj,�P�%�W��Y�8��r:H+p�H����2���o��m\ �|��'�8_���A�'�Ȫ#Ƽg=c>ܜ
^@O��ˋ���d2����O���|wٿ��|&���{�YX\�R-�A1ܦAmز�2�jl7��j��g�d�Mg+~��(G��p����1>U5�����?�}`&�e�X��N8���9���������������P�#(Y�sgU���"{���7��n�����ӡ�ll1�얮,y6ʎ��'��v�`b=����j\���q�G?���B�#|a@�>N��R�#oKy�X�M��=:@j��5������W9��=����e�"΅e��趎�a O��o�G>\��޽xz�n�?}��9or��pO�+�[����sq���x��7l�{ۻq�}�)%>]������{o���K9jBe�>~�,���}�fl�B�������%�����X^��[ڔ~A;Jկڜ�N� ֋���o���s2(���<���Qن��6��>p�`�;��*��Cg�@���ϟ<񦽻�ǆ���1���P���t���[q�����W���8�w���~���7q��?{���vqݑi:ګ+џ�m�Ă��7ވ���޿�1�Si;�QJ��$:H�������_J���� �ӎ��
����q�d��N����9���y����=�<��[q�?��Ç�_��f>}�(����~�8z{x�q�~E��Ǳ���9�����������9�}�3u:������n������O�z<"��I'�(��\�Uz���-k�e��'^���q�s�({�O=p�mL���a��a�o�-�1���ƶ/�L�I�ɞ���l�p��n��(�>b�a
����;Rc(�� ��$(�� p4-+�Wp��<��{���ޠ�����C˲��t�.�n �dH�iӒQq��^HW� �>��r�Gwd��\�1�
&�m�7�La/>���ӕ.K���o��O�����р�K��P��i�,�s���P5y.3��8:B��&���34�	�+)Q�zDCg����6�A|uxwJa��P�f���f�C�zp�&�C��/�hy�s�	݊S)ud���`؍99a��۱{���3��7�֕);pS/�+��*��$+]C�[�-M�+����/V�z�u���7n�ͪ�ܓ�`%�N������+?i~v���b�c��w;��AՃn�շ�>��4_c
�<;��C�8���$+��fON؃�����>��n���P���q$�!���k�v�B���;v��e7��[vZ���a��x.�Ԅ�����b����ɧq������>z;���'�;>�$1��i���`�q��t-Є~�9�o��Hz��h���e���� ����8bS`�Hr�7۳������)�g�楏�l���{r�����W3�7ף��Kr�^���_|O�h�؍9X{�;q���ؒw�����G��훷���-;<�#vxxǪ��nŔh]|�m?S�q��d��=��Y-��8��!�������<i���n|�NesBS���m �Y��|��N��[R��:���a7�_x<��W5��ljA㙟�:������P����(�|ON�7���{�������$E�/tT���Z\�����X���8���sa->���:�ua��F��)�8M8.�[w�ǎ�Pis����$��_s�>���� �1
<�d�����v�i0T�,+����x��an/���w���&
 N�df-���l#ƾ�����~�q*�Q9�? �f,���icc��f3�p��I�e^Q�B���������ӟ�ʆ7d�V@��N�Ƕ��6M9l8Ӳ^V��<[�|�T���κ��ۥ�6Ϗ�+����'A��/���w��;a#C�3���cM>4�p�����6a˫ �212��Ni�0���.�8�L�+�P9�74��*0pq�p'Tx�r��&O:Z�L�:��7�(�|���'�������*�2�5�$����,|Ғ��2���5�N�Ny�inu����}]�k"]Xh�٬x��g7�hy�r���R#��׃�d��<��� V��AL_���%�.�N���Y/�Nz�0��΢OOmN��I
Ӡ�?����!A���|���ѩ�)��S+����dj�Ǝp�m�I_�oi��e=���u�:�C�g�x�����ut';{�6;�����b�����>���{?V����{r`;lɠ�O�����Ə?�����,�uѱ��7q��&�?�<�=�`�[�}^���ړ����=d7����X��>���J��RM����hd�h\�QMN�|L�X��.�X���	'�T�e~cO:��ؗ��Q�SQfK.�ߓ�{�������ۉ���xq���T��bz��M.ą+���#9핕���{1\^��X�{r���0T���;�{��a'���x���g0��ťX�r-V/\��C92�O�A��s��/�4��`�S':b-�ϑ���|�"\.�(�*F�^^x0q�-A��-?�*yk	�U�{Z�-�m���@y�(o��^���G�����!^|�e>�g�C�ŉ�M�i���rt�x3.�����_��[oǌ2V�x��4Ҿ���Δ�ER0V0�`#�	�e����̡p�� ǑƩ⇜��1��F����y'�ʣ��τ);M�8�l��-m�M&�#��|Tv��9���Ah;��#�r��O��C�o�=.��nʫP����d�� vl��� �C£�)G�1�sxq^S�8�|ؓ�6��z�J_&��\��*�e��8r�N��yݔ�#�0b�O|�!\Hq����j�T��+@{T_��_+h����ˆ�;������?��%��t~1:����,O��UuM�����l����b�߭��dY��G `3�2r�"����)*�MU�E���5����t�$�Ь � >����J�����T�C��\{ݣX`����q�����[ў�� �`�%'@���)��y<���O�����*9V�f�=�֛���_č_�"b]�<WW�!�B�u���bjq9f6�Ō&T���~e_�KGW��N��4O����^mE�	9u��$C�(
���Ҳ�EQ:AnOpD���ì�2���rGv����c�����r���W��F����?}?Z��}�A<��xr�n��M������kqU:��j���ob�Ӊ��a����Xz���m$>�dGK�7[�0���s��P=?��?�Q�/�~�Ճ�tְ5ٙob�h�:���� �J�+kl$�k�������|�Q��$7��\��-ɮ�����8d�Z��>������/_�o��v,γq���ȶ��1ݚ��㣸~�z���`�м���=|��ݏ�>��+d�ɹ�ʍq�ڕ���~��-<��@&	���t�]�'���ȗYD�x��Q��|$�=ۈ����Ln9Q��%i8^��ׅN�Qw�͊�)��"���{/>�2���*N܏��s�B7��H��rZN�ڱ��s/�ʇ?���F�=����TN�$3�\D����^���:�g��N#_m�<o��\���+�s�Z�T��J��8�.6G}K:�a�6  ��IDAT��v�mK�1�gZ�*q�t� S8���
zu=�>��`�WsB�M򗫂8o|(��L�&\���)��s4?�A;��\5T�����>� ĩ:���N�̵�<I�t����&�8c���M#?8M����&��?鶹hQ\�h.ae�c�,����՚�*.����g���o�g����J����3N�U�������dl���A#...ڀ0�rVҨrb!���g�,~t`p �vuP�+��4�>���s�<(�H����(�z�˷ �)�K�o�W+(�4�L��� ��m�p9z�<�(t��O�Y�_b8y�N�u('S��P~��tig?��<������x���1�3a3�弜���XX]�s��cY�m�F9:����fc��%�ڇ����7TvV��sj9�$s��q�x�$=y�j��~�a��+�r[4��b��a�38����%:�;=Ml���W2�󚺮`�4qO(Jҙ�E{P��n�D6m�w�H��l)oM8�������z3��W���d~����[��>�"�����>|���rh;~���ۯ�e9Q��mol����8�ٱ�ĭ&���ט@qphG��=Ȋ��\�ލ���[�֯�!�W�ƱX�-Ne�̛�ހ��3�r�2#HJ�S��u)=/p�@�K�x��29��������^����}�qƨ��/�9�	�{��^7�r�ݜ atkg+���)+���w�¹� ������?��Ob��9���g_��?�(n޾�.��e���Z�����!'D�҇���2l|ɤ�]P��G�L)�}S�ṏ(7W��LB�H����.M~�ES<��Qt�c��d�l�K>4�ƽ?�!˱�}�~��lg5Av�;��i�ݼ��z'���Ǳ��;1�*�S�|kR60-��A�m{xP?����_���c���P��?z�/��M�)�!X	�n|����o�a�,��G�d����4��)��.�LD�� ഋ��K:/��T�<��������/��/ٕ�n�82��j�(����;3JC����Fٚr�e�q�'/�'Ȯ��nr���X<�>�m~��H�+�s�N�OҶ,j/�N�8^Ԑ�Iڰ/:��6����z����z[�͝x�w2�K���Sτaw�ގ-MNT������_u�jT��L��_?h�d��:�
��A:��7�3�������<��%z�� ڤ[e�^�e��$ẲN�o�C��AŃ�p�_�ns�c��w�:��O�#���>HE�9s܏���������F�);H�.��w߈��_�����
�M���B��q-�k����]_� 2@Ϳ�ۏC9u�>�,�I<e��oo������݋6W|�{as3���G8\�s��I��gC�ǒ� Ӹ�O�
F��X� ��w::R��9������S�+��r,�����b�ZS�y�j��ßǢ&Ż_���2v�?��&ө^?�j�9]���;���E>��d˷z�|�̈́�@�A�%�����H���{�\�N����Ltt�ʂ��%nũŹ�XL���6�<�>���J#M;�đҍ��UVxJsX�PT+\�{���ჸs�V<�8��?�}6Y=8��ɷ@�vwc[N��g��ѣ��b�mw Gzn�Tԭ���ʘ �>}��݋�Дc�_������O?�4��m�,�/��?�~��x,'~�� ��r5@��|����``�0_�6��n,�dn�Xd���}$'�W�0�i��5D�h0t�g�����#i��A�H���N�l�ż��[o��eEѺr5���ø��/c��Ee)#��S�6T}�������1%���
t�V�E:��% ;�X^�$3N:4tI <t�~
2/q��%���8/�C�d|�/�渄͚NC �K��x
���� �@��P���2:���^���h�<3m�LO�\o�����SLU��
ֳ�$=��ǳZn�~ѿ�M��t!`�4-�%/�2�0>�/���`�����i+�N���܄�f�^���hu{�����x����T00��6�Sz�bHc�4�ȸmDJw�>EHjb�iU�:U֝PyU����{f�QZݎ�6h���[� �����^�j\5-:V]a��@k<g8��eF@zɚ���RJ~�D�~<pk���J�.�|]��w������/���O�T�Ī��׮���ϟ���a|�����/���17���s1{�B���q�G�E����Ɠ/�����Xt�x_�� 4���b��;�7n������׮Ǳ�u�[r����V{��*,�_k`A�/lH���F����
@�=�\r6�o�J�g@<��c�I���i�Cȷ2���������\X��+�����x�����7�FLN'�3��%������v<6����\-��lo��R��	�[�}V����X�v�{�Ņ~��u?�?��3��m^����T�C�@�pv�F�I<�����ζ%<�ö#|kgkK���x�BN��a��R�s�Sq4�x�{�ɀ�y��M�yc�}�� �8��Ҿs�c2���O�VȰɣn7����6%����?�������������۲㈥�u׃<��I�~�>l����[T�t�x�vnt�-�𪌀[V<�N���)�{BS;R�d�)4Gap&���� ��xˮ�������ًx�ۏ����S�+���z1}�b����_�2�\�����]/����R{�3��J��|��p�`%o������t$:yKR6���C�N�|ƏԉS}�Zi� //��0։v���AT;+�s�)�f����@� &�*�|$.P�\���{�Vļj��|a�����$��Y�s�;��\��qy8�.΁�u��e����M�6Y�s[�=Y=�tpY	9Ē�+�f7�+��k���H�������o�#���o#k���
S+a��u�[ߓ�޿W���-ނ��pq^�P�Ё^m|�P�4��;�\����Ǩ����]����R���ܱ�de~��3 t���*�NZ�r��i���HK:���~�����)nʕ|տz��r �J#����gD(��L�\�ȁx��Q<~��{3�#���e\��4P����˸���1��5i3Q�E�[?�A\�]�����q��9(<�~����ݘ>�#��-YϤ�ɽȎ�K�v��.�Zr��<��0'�v���<�Lنh��� �3��k�Q
4(����t������O����v,��z��O�������O���Q�:��g���Mm�Jc3ט���ι}�'V��ϩH6�f��C9"�8-r~�77b��kq�?�7~��Z^�&�9��	���A��B��iʉ��㈐��> ���h��m�3��׽;���/?���Ǒ�q>6��f��!�\N��U�c�a��t�u���k뫱y~S�u?ƞP|"���9��Y�9������8w�\,K��9od˷"�)w�݋���q����_�wމ���W/_��?��:��EN"s�3�3d�����Cb�/��-v�����ԸS8p��=?��8��ob�UV�x]tY�*>�gŘIp^6n���'���ub���R����Sd������ď���W/GGvs���Gu���h��N��g�a�T��EU��E�����V��țzH~U��3�'���8�F��S�@>6��U��)�W�_<�-N�ɇ��m��W9��dq���6c��QP:�αɴ��a<�]��6�s�H> h�ؘ���8Gg�dR'�P�6�(6�'�BoBp�#�GA�-�\�#��H�w���3tG9ҳf��<蓮�Z�CE��؏��ƣO�Z����6�L�k����WC�qww'nݾ�+�l���4�F�`H:���O�lJN4�d�;�i��0Р�SC�	���=�V��t͗��z��C��)�\EC?�)Y�����ƃ��nP�`ޕt*h���j ���e�|�]%g�����k7OLt@׭#�ݣ�x��o��N��>������g����_������h����4�j�`2�z�,~u;���8���;�/h��$���)9b�`_�~t���5���XXߐ��AL�F6��p�X!����3+�"��B�o�&�ǉ݁I�t�v)=5G埴WϞ���ܔ���Ho�*e œ[wb���8�-g���-p��q���a �<��Ў�͵ظr)V�t������-G�L�5i)��Ĝ��ƥ�ލ�|k��~;by9:B:�·R�U��VC���U�l�1�G	]�lA�H;n&y�'���on3ޔc�ŧ���"�=}b[�6xޫ%="'|�KSv�VV����bS�պ�GsQv����¼�,9c��f)���j\⫊C�g�܋�{:��a�K ^�<|(�����o��4n����Ac��V
���xH�86@�����T��s�b<H�U_J�ydՂ7�?�#��fr����L~t�})OS���*m{Џ��x�׿����ױx�b��	e�wF}b�L��<�7���jW��6���v��O=�odŲ�c�z�U})��s�&�F���:ih��㩷�G�?~�/�JD:N���'�\lV9�~9N�O�3��sN[Y��1e�\y~�_?���2��3g�t5�3�p���t��)��喸e���w�)�oy�<@�����7���^�s�{��S�l�̴���,j�.�%-��<�
8@�|�vN}z�_�����V��.�t�A���p�Z�{�UC�Q��W_}{��j|��*�؄Qg�x��<���*K�sa��44c> �5M��$_.�䧱7�4��<����Q���B�s�iC�d˸���Ӥ�s��~�K*su�5�.������<@��bU�/?�E\�tQN��x|�v<��Vt>�V��5��̼���x�<�νع�ط!�ԑg��ȅ��&{nC��'�~�f��j����G_W�|�pjiY�d[��Q��B�U1����C�&>ҙ:�l���J�l%u����<��j�1l��^����"�5�|>8���il�y����6�d�[���V��.�¥sq��ո|�j�[ߌ����z�<zG1�v��6çn����݌���r�n��G������kޠ��)���3���ᣏ�F�%�d��`5�&��1'.��q�?���޽���?Ɲo�����\�{� �7a�$�1A����\ˎ�2��ˑ���m���%�-�tA�v�s?ؘ���Q��&�#9��;V��\WVWbM�y�Ϋ
krHW�W���6wO�_���Oǽ���
����{~S�7:y����$e����=�'A��ڼQ�u������e��U��"��#xI�8bv��(�c��o^m�y�J,_�����_�,V��Xe��[N̞��mV+���Ce;(>�F}��5�YF��M�읤���2�fh��!9�U��"7i�G��#�rLJ:�ȋ�s����e�E�H�_|��?��9�h�^�^&-���1��r��wK([|�����C�s�+�*K��<�|�/\tctf���z��N�c��j�����$��ަ�c֕���b�.C��I�<�@]%�_3|���I�h?��GJ��β�
��+�H�VY��d#��*��W��a�:��_���U�8���>���y�IY�*A����c`R�N��D9�p��诉��,�Q=�a����z�WhX��� ��FM�D �z�_�׍�^W\j�_l��kW�ƕ+q���>�$�U�3�;!�6�#�
���o��I�˺�_�nE���M㹣YՠA�GASN1t�{g�qԚ��r).\��?w��� zB�C�*�I��'�qdbh�f��2�MU(�Tv�*C/0���Ωړ�;܂E�a��7�=�no 'SvM�/����_����q��7�q\M��l;��I=�;�|&
8W]��:>�ɩ�*l��7};�duɴY�:ũW�N�XRx����>�ˇƑyJ����@#'���n�s|蕥o��:n�]B˼(C���پyވ���ۯ�R5?�������l�/`�&�䜱jppx;��N?�����cJz�u�~<���lO
<����n�s�g�A�ܿ{7����&�C����;qK��|�;A��*�̹y3�M�_��F_ }�:k _9��H�V9�s�#o���CtM�y�{�E6϶+l�1%n\�W�z3N�])ǫ/d0n�s���0(©�G�/~F� ���c# ����82��S��;��f�Q�C8�<���,��F��Kݤ��9dZ�.+L:�͓�#B���r��;��g��<q�y��V^���C�E�'~���L X��S�����Q��J��a�!�/M���P�M9��I2��E9�=ҙot�#�$�8�y+�V� �^x:��.����Mu�9��L��C�� �3��c����S�L��I������3a4��nݺ)C��a�eHj�l�<3а
��9���ƃ�wʸ�$�G�z6�ҀI����:���o< S�~��u��2�Pj:CCW��:M�)��r�ϐiY�8G5�tJƎ��p��dh�O ��I
�kO�3��^�i2\֤zzt[w���O?��{����X~��4��L������2�h2�� 5s��fx�K��������/ke)�/߈s��}7���ů��N�fJ�V̙��d\���V �� 0A wB�3`/��� A��=�юԭ,+m����ǂ&�5��m�g{����{�ܺ?M���~7~�~l^�S)g`k7�~}+�?x��n�}9��`����Y��h_�������[����f�,-� �O��o���Ӂ��Y��%3OpK.��Ii,i9Q((}(���n��o������n݊����W;�;�*J��8^l�Ж�y{q�+a��t��Y1Ʉ#֓Cu,�y��Il��Ƌ�/boo�[Hxլ+����*���i���Q��l���h��Q��öU�,gpT��f�r����Nl�i��7o�ln�����M�� ~�1B��M�@��L�<���Lj�X��*c0�BNf����w�?qq����i��f�K�$��Z�y�����[�<�G��:���Rp&��	9��Q���<�I��L��k�?�;����Z����11��8}�t_蒢lt8����'�cС�t���j�3	�;��A;y��2�����v6*G �l�_^\��o��)K3GP!���"$�n�'���My�iһ�$�42��&>|e].K^���YP����C?�+�g�y�
�/��}O��j��ݝ���x4zu��a�(���L62�E�&��5i�M�0�+Z#���M����z��I��	<�4F���2�F�:Is|�������q2��Kz��4�<����*~��Χ�諯� /T[	-��԰g�������1�#l{ߟ��[G0��iB�9��ɚ�v������DX���5yk1�f��qX�9k������x��|��|�������Ϥ���!�÷אA|����X���:4�(������P�x��.����m���J-;��ߒd�B��z��%��˯y�Գ�Ÿ�ޛ��~o��=fG�{��?��_~��P�Ĕ&UoQ���),��ٹ���˟ƕ��8�׮Ɖ�v�7���rJXL�f�Ɖ<��"�Ǖ�&d�q�O��[�<�Ęjc��铧q��W����k<}�8֖�cqn�_`%�ېl9ǭGMr���ژI�CMZ<�tt��9�
6�y��C9E=���q�qY��f��6$oD�'��J7��m���Ǐ�7�4ซwUu��r�t��r�x���������?>�L�vpu��|\����*9�+����LG�QܧJ�O�ߡ�XJ�"-iA;ml����Q���ʰM�)�U+��f8ߧ%�1��nk�R7~ك� ;[�?U)�t_�����+���<�z��^�n:��H 2��q7�H9�ӌ��^T�pr�I}7m�P~M���&�1��]�݂tZX*~����H^�k��;K�K=�@<���d�^�a�_%#G�0�r��U�뒼�I%��0��kB�'xN���t]��N3)�{2k�OB!?��v1e�*���L�"���J�C.|�D�e�L��gp�Z@0���^��?m�+E���?������x�>ԍ���I�i�9�,�d��*&��4��y�&�L+��H�� F쇜<@T��Q����`�^��N��x�9�,�3$j�G9��ߘ�WOr�r���4����:����(S�%R$=�7yS�&��/n��98��dЍ��8N�>��?~��>�����u2�q�7���s&G�o)��,�:t�7����Dqp��ޡ�fˇ3y}]U}�0�q���q��wb����]M�gK+����r��ж�05?�b��I�!��*O�>J�9���#�M�faG	C^8`{	ޚ�����Ԭ��/����b�n�It��ŗ�ݚ=�%V&����W_��>�]>��ݮ_�X�I&n�,�cOf5w�rܐ����~�j`�a���y9�<t?{�
X��t�	��s�lR��$���^��=���������8~���q��"V䀭,.{�I�I�v�o��l����l��~�+��o�.�:-�ŋ|�ve��J4��I�S:K��1W�na�?y����ʗ�m��|+ӧ�Su���q��e�ϳe����LKr��q��s��xtO�>/ӱ����\�S�U�q\U|c�\ll\�V[Nf{NN��h�&Ydæ�����Ls���qI=";��cAfdO�ȉӧ��*$��4P�ݩ��Z\F���4q#z��䕝
����&���l�r����ӄ�����G�<�I]�L0�U_A'��"20���}�G�'W� �kl'��E��Ȏ����ǭAH�o�?x�)gn��'хwꘕ~Ŋ/�j�<�N~�m�<*���<�Ф>�b���J�&('�j_߂�9sX�Bp{�4�`�o�d�[�B:JO����'�:J]�Wu#�&}��5��я��j)O���������<��2�YO֛cj����=p�h0��pCj���lk�E��7�ͯWϷ��pD�g�t�~�ah 8��L|�^U����N�>0�I�+��'���ʠ����
D�®��
t"ҨÃdӉ=Q6<=��W�9�tҰ+���CPEߴ\_A҃ϺҬ�LgF�#�dH'D:�?#��~?�<X��]9b_��������a'O�LyC�����Abu!�/lh�[��0�3dG�_x���&jx�9#���'S�р:s�b\��q�G���;����F
�+��	�F��OzA�̴L'��� ��kND*��=�5��˥}"��;�=�`�l;ǚc�sՋa�����ډ�Ͽ��/���;���.�r_lO!��r뭯���q�?��>�EL���-�dL�1uV:��uC nC��?m�N�B��E��?����~�,�������/�sȅЬj��@�N � ����lV� ���T9�Է0ߎk6�Éu��L
<c�dK?b2�s��6V�X噕#�۔��A?V����rlm�*�Fޚl�há������|�Ď�y>���5�����a���kq���^�s�.��t$9��Ф�S��z���>��L�?����I��}�|q�����I�O�/� �V����/�g}��̣�wl��y�O�r�_�D� �M08�~)�+���Z�j��-jhC�(��������1�8�qN8�sL��\|�R.�U�u&9tZ�l�]Ǖ^� ��6�sх'A��6�T�sV�l[d�/�ĭw��@�g�^�)(~88�M��N����S�U:Y�u���L;���<~��#a��ϱ�l-��o�R߻�(f<@Wن/��]@u�_u�����v$E�i#������Ç�zh�7�#�@00�&��F����I�@d�1q8�;&90X8��Ǳ�$���ɺ��|1`�	H����Ѥ�2x�� �tB�/4i	�ʺ�n�UG�����$�w�����X_[�����"��q ��K�b��k����q��7�7_�e����g���I��i��.��o�>h��[H7��e9`7~��|�����:=��A����7�R:j(R:��3�S_����
Q�+e}���{���im�y��8�0-BO�q���_����t&ގw��٭[��˯���ocF��	�A����:X]�����֯?�7���܈cv��⃺$�R�ｼ�4�a�͟�R6��O ��5'C�1�h������7����΋���3���BQ�9�p{`gzdR�\x�C|�(�9o��ɉ�H��~r=�����>���Z�ωu�̑��?>�3c;�;�����U���q�ʡ=:<��j�A��6�ެUΜl��׸��߸���WQ�^�k8�ܚ�_d�ʊ� �h�I�INth��o�@��Ɍ4�&Ǉ��u��M�h��i$�G�^٪|J�xc��Gy��9.q�S�Ν�m�c�H'
�5$��O�3��l��Q�S`��1�&��Ǒ*�7�P�p��/~��H���w8 ��Pu:��QEKǖ<�Y6�]G�!O91֭ �/e�8D%�a�V��K ���H�2��B�M�ZGp	����&� �;&��x����i��ëYN��v�P��9�?ҲݒG���ߤm�@�GP�U�k����9�v_W�|�h�W��Ih�ڐiXcp�~6:a��F��|:]f�IeL:N��R=�R�����D�t�LfACWR�V�!�R�(ޤ���"�5u�hCqN�����1O��d5�R�Ҿj�_O�Q�r�EZRЋ��uv�|7��1w�|\�ླྀ��w��߉�
+�q����:^ܾ��}9�6���hU����ސ�&���/~�r�f���lVe/߈��+!�+ݠ,r�{ ��Q]^�C�/���W�f=[/d8;A�º��2�{�t�L��4�JW�R9���A�>~��Î����+��j#z�9[����Jl~�n��˟J�D[N��rfx [uC� ��نe��A	��/��k�r��|P���Q|�������8~��9o���5�j�*�o/�3��^� ������m �G��<F���<�,Ⱦx��~{r~�{�������Ȋ'��$ ��1�91��6	�g��z�2'�(��M{B��~��ǄI����$���[^ZqH��q�iK�q�Q;���)1oCe�W`��tlT�����d�t�ϕ���£��ݚ�"�@�N�9fT�ğ1�f�W���XG���{�^)Q��GuV�OZ�̄�,oFII=�P'�&�ꡭR��W���Te'��g:ē?�9-*������Jnx��C�7vd�\\�Nt���\:Бsud����$%铼����~����+@>���N�9u'�
	��e��<�O��Jϱs��L��I������'�*#Z&񊯿V�^�����oݺ��>���p��oh�
��*��M«�eL5@�:0�����6X3pT�>�V)R�Ń�i*p0����8�/��&@���@�m��¦��
��=����#����My�w}MXNf������^{-��_�+?z?�|�v\|�߀��f|�������$8�I���U�����1�EM��݈����v�^�'����#���5v�g����rJ�I0m�!��2)_#��RrbAo�/-���v�t�4re)����f�*9`l�0-x�����ã8>8��� ?/���f���Gq�?�3�~�t�Q}��ਛUH��?����ΒǦ��V�{n&=V�(��xfuM)lC������8�ct��f,-ʡi�_�ղQ.�d�
g�<�۹�	�*�9��lO���ɒ�����EY�������G��<[I���DA�[S��GvP���A��6	�N�G1��	ת���?�g������u���)Ռ��~��VL�dzu����f;hҠz��O'^�z)ñd�6K ��!�y�/D��D�cGڍ:�0CP�S�+�̤�Q	�S���9�~R�����XY�q�)|�f�̶(���蠜��}C[@��)�:G��(�z�>�_9�TH��sn�[�nN�W�2�lW��|.B����nzU��T�Z���L%�d��=�[Δ�X����I;KY�6+�e����,C=9~I�����
�������$_��u�0�����ͯ�FG��7�;�x�,pG����<I��*K�۱��e��j�A��)����������y�$G gcz��p~S�N�Ԕ�����@H
��O^��JH����g �t��ڒi<����G�٤��RCMh��q:��b̝?+�.��ƚ7j�{�(n�����ǟEG���a�t���Y�XӐc�U����7ߌ�~7~�+o���SѕVSv��r����9�2 >��Yw�){! cM>ЬvO]$��v9��c	e�� �[�"'{�Q��d^_Y�ե��w�Py��;Y���7߈K?� ���'���k��`�;��]њ>S]����(���N.��,?�N��L:8`hc���W_|����]���\�ܶ��N�9p�����D^j�zȇs�s���Bxa�[U����ˀu�s�����.���#�F��/�,-/�>e�5�)��M������~��Almm[�Ņ%ORܪD�M��I_bE�@��{w�nll�B���e\��K{c[��quч?�$�L��|�Z�H��$�J@:y��d{�~��ӓ��)�M\x�04���}$�i�H�S�fXD�	{K|��A�<^g:���x��I��/ә��s�θO&[�h�LE]&�}s:څq uд�B���9Qdv(Y/�e �C9��6�2����}�O�&�²/�l/M��B���tL9��5��y�q���:϶�z(�cʐt����6M���h��E'��$^��.�������J�{��~B���5V�@
TCЈN�D���I��i�*���':���8(�4M�Aњ���x�.GOD:�F9e�+����rY�S�(\�YF�� yd�/�v�x�N8Y���`J񪜎�����'�&���>Wur�-��u�i3Q@�j��6�ˍ���� ă����?|��q޽�ÓXP�N�(N����C?Q���ߏ����/?���s��ɓ3Oh�p,��[n՗�@���ޜo� V}�ڃ��� KN�A�i�n�h305�ה��z�:����/�p�9��p\X�m�-�`�$�llně���t��X~�g�g�p���IżA*�i`�e�/�+~��l�R���#oŁ�	|y	��o��������&�>z�m���y]鶐[�"F�qT�C{�S2�#��g��zD��_pq����@u#���Bꉠ��Oh�[/^�����}�3V���//�E �ͭH߾�M�A�%��[ԇ� ��xxx`�	�V*��}6�7�ٳ�q��x��>4���gl��%2��,�s������g�e�����Z����"�d�D��;�36f�������eڦoUWu��E2�d���{9��:|��d2�#��>8��p8�/,,,�9���c�+xN�C�,�	����q�O���5uO���IZ
����!�ɏA���>���VxFA�'}I�@y9���+yp]�#ڌ>�At?�?�V�׊3}b�T|�ܲl�%k�c���s�6t�s`z��T]x��,��o�N���U����_+��B��L�H�Z�Y�ͧ�Z\�V��V�<%����U\�ِ^㏓�XZZƑF�����|'���A��i�I���w�
�S���<o��4�hL_�}o��&=z���� �I/`�Q.��S�]��@�+���A�8O�Eg'mK��(�ˣ+�69������3}ьt��J1�쬩��O����1]\�@��9�)���JU���!ۄ� ȕ��L�׬=t��9X��ub�᣸�������b���X��5�����xT��X쎎���R\|�����S���'d��.��n?���ec7P�ўx��Q�~�#�oB�� x�v�Jq���H�* ��J����.p�\����q��c���B�Iɸ:����g���ozlHܾ���G�Gh�?���5��4�Øx�笃�p(�<
ϟ*�~�A���'�k������N,-Ƭ��PES����~]�'���`��!�!Q%`�����Wݠ��WV�X��x�q-����)ǲ�_y��W�����a@Ꚇd�q�t�<ȁ��y)�I�V܎1?���د��;�����]�>�?lܿ�7�L68��7⨟�R�%w���~���Cx)�6��{
&7��7-�t�=���D��S�&PJ�5ˡl���}�Y�y�D�"��������a��w��d0*d��WU��l;��¼8?��[��NP5������oң,MGL��V/9�C_��pE%ˤ���IPx6 �O~%9���!��`�G�T�z�X�X���r����YmC���� B��%�y#�L��`=T�+L�A��9دw9t�5c�����&��M���6p���*�_F�0�ty��<o��^	c����~�M�42�EA�{��R�Gv72����kx5�o���
o ������sOQ_�*M�z��AQhU[��M���RH�,�f��ؖ�<6|��f�~E�R��M
���.�DX�%i�A�O���R_O6��հ
�9ty��5yu5������9ڏջwbge�2�1��V��Q9�'Nǹ�ގ~��8��[�ϣ�Ξ�1Σ�'�F��Q~�B�^�3�>�O�g�5�Ps���{�GE����\IB9�~�S������r0dLr�,�);�҅�Qs�A��r���Z8w6�O�� �%�aL?Û&e�)�,���r~��Ay�L,��_!�~����n'֞���/��_��?���\�N��Z��@���$�Yw��r">�+ILƬ�Q�pޘW��l$��EڼaH�"������e�ф.RV�ыw�	�Ȯ���`�ea��ʥ��>�f5���g��nJ�>�H�S��-+`�.��ǧԉ�]�����_��Ќ�3MZ���?�����|[�8K�6z��ܖ�F�O�}�B��c]2�c�\a���_�?��>~~�<�#���K)��;Ty��6�l��1\��`d�#Z^-٢S�9��cPi��vzZ��~ʄ�e%<��p�� >d{a]�j��o�ڃ�u���/=[iYF�e:�«�&~"L[zȷ��:�1�9����ß��/�h�ﳴ��x0>�̱W�K���98�&���Yb���2��A��O�����v���[a�%T�W�W~+� �]���\_�!�Ox��6ߕ����z�!j��c.۪��̇#��R���'43�h��+e⅛�g���rQ�������H9� ��uU��u#.;)/��\N�%#]�?銠콣�����&䡘�����~����Q��<g�|3.|��'Ϟ���	sD*�ΨFptZ|�,焜�ԉA��d!�̿ �M?��Y`�: a�Qʐ����i�����Y���*O�Jʨ�%�ځ�rÚ8F5�c����	|�]��$?m+�ːe�UY"GZ����v&`H�O�g����ݾyӫ`��v��IM�≉Bdx���*Z^�wQ�q�'|�0�(�r1��1�����C���8�k2�X�pF�L��� N�7M�C:���ŵ�t�.!e�	��V�l��hA�p;��~��ǥ���0d�#M���G�,yK{qiɆ�WZė��@T�����#_|M}���/9�����Fdbn[9p�K"�ϰ�t����4�F3�M���<�g>�Y��c\qC�Y��z�I�%���ܩ��������xʲ�O[U�k��F[>�~�O�3}��懇�Y�@�p}���rh0m���;��0������+�p)�x#��>����?}H闿�!���DOg�sM�E;�?��p�����8xC,�f\��
������cc�g�}�;�P��r0/�%�{�T�X^�O��RX�p��A�U�)\]��� $�@��s�[<q��Dr�2&i�0������\ɀk�e�����h9��MX�8!�ǭl���)H�r�1��	O��v�H�i">��!9MlݽX�،�����r%ξ�f�|��8���1q�L��HNƛ2磦a�e�(�}筁+�rTJ�t�~0�8�)�QD�Rά�X7�ǿV�A�����	�A�&B�,J��n%�5����EOze7ڊ��;m+ls)�ڬ�#�iB2Ax�����f�@�Lzm^�q��B@�ZPq<&z��q��W���?�$.�?�u�*�d ����VV���Y��I5'�\�gV��eRT.��at��Ĉɟ2{�;�i�������� ^{���\�W��(Y�j\؊��͸w��O�����+�96�G�y�~���[ȣS'����TY!^��_>{��%�Q8�1�O��ĉ1�ɇI�#��R����E�n\��dD�ȱ\�+/L氇K'm��W�
�I+]r�P�u�x������`|r]]�j ��8ϤY_�:�WK4�^��'�;Ɨi���F
��/�P>z�O~ʢ��S�}I>I�/g��2�����O>�d���?�_U����e�N�f����ӈ�my7�|�'D��?��*;�_�����f�U��J����͟4���p��G���4< Rx�Sqy���)�H��)g�V��S<������������{�Nܻw׃��3��},:�EY�QZc��F���}�������<WP��g->�Xq��5`�6�*ݭ�ӵ������G�G�Hi����O�1;�� $�?$�
��ʘ�zb IR.�Q��c��xO�F�8�<��g�NŪ��M\��y'μ�N,��z�8��YU���I�X����C7UU��ruI�\ׇ*�#���� ˲Q>�!��4���,������C�mɏr	�������ȇ����#wV�;�ѠǷ��G��e�5�<�R�'��Ȑ'[��rNk~�ߓ4����_�˿�ǿ�m�NOřS��P��B%p��1��|��*�Ɇ�Ƽa]i|����������BG����7�dа�c��ٹ8q�D��/~�7���F\����ܵ_�^���a����w���Ũn�8�k}mC2A�*]��&�mP����޹����H�O$����:��71��%� ��0�4#������%�����K���W��rI>R7́��a]C��֏����@�+��*���h;��٧�B��&o��K�L�5y��R�c��|v��¢���'�o��š�6�
�xږ��7<1�s̡xV���,��'��,�Q�'���+^z�a�dL�4�o����L�y����˱\R�.�y[Z��P{�H7�J�x��0�iNS|ѯ�H�.�V\�#�Z���K�@�e=-�:��h�� @���i�*�R �S?��2~(?}�~̛�)�|^||~��O����nF���[����:G�_�/dokp���}J���hUu��H�FgP��̓5��t~��8�k���2 ��ф��E��L��x�|�ݼ��'�N������AJq݃� ��A���"]eP
4P���	�1����Z�*B��c�ܗ�?'���[�"�ӳ\ck���1Md��6�g�T'�?�ĸ��������Oӧ�c_���$#Mx{5���:du���`s��Nw�^U�@ �έ���=G�a§�݆��2=%�މGm�k��Rn-���!��f�����<%�Թ���ަ99�������|��q��BNߐ���L��ɫfr�N�S�+F�����ƃ۷�����|�{n6�磳�k\�p$E��:�A-�W���G�s�s~t�i����Ͼ�hs��~��u����Ϝ�5�8gZ>�B��n$�:u���#y��ۤ�ϟ�s��E�Ӊ�?�8���!n޼iy�$@����N��Jy<2�w�q�<O&���77��6���ɝs��=x�^z5~���k�9��L��i���>r��(7���(z�x�_*ŏ�o��2��)�kʶ��"<��8�(ʕ�}�M�Q9�['9^�� �����+{rt�<.B��ӱ�V7���r*�$ԥc���@��ؐ�ܿ;�jO�S�ўt�쥫q���V_�hR�*�ߚ�z��]S�{���	� ���7��)�Z�����xڬ1n\��7�6������>��<� �cs>�Q��� ]t�p��}cI�/9cW�7C������\~ӉjˢO<~���h�s�U��X����=?�@OK{Fb�/m��̹�7p�n�^y�^��������?��0��ӓBi"������}f&O�F)Q'*�DbEUãP�S��cr嚯gc���!���j%E"�0���<M�u%��~͖�(I+ynE�!�=�e�S��!�ɀ��!<�Q��4�e e�OqТ���=bO�b� �z�m�z� ʶɁ�NG���b�e�b��(]�Ƃڄ�wV&�\����c�1"Ŀȱ� ?�[cJ�ٖ�~��r\��M�G~x���AMGl�(�q��	���H��r��8�c$�<�_n����������[v���8���聃��Ы8�8 :�y<u�@�<J���l�ɏ>�?z�}�������Ř�S>j����Z}%�o5*����c�b�d�eR���	�1g>�OeX�9�~��\�'����6ܘ�S��3�<u�߆<{�l��g?�k/^�ߪ��?�)�ݽ�w�ٌ�'�Kۏ�N٘���'�?L�� ��M�$�Cݺ[;q y�"s�G+kq��J�_�����|��X�!�J���Xl�p���h١D��.Y�\�d"?��!�_�����s��q*-@^�X���r���C�1	�St��4>&lꍼx�?94�|L�H�$��j��ё!�����qՀ�ǒ�ڃ{����X��1��A������^t�&boj&fN����F̽�rL^�;�	ubXTvT.�)nK�ݞ�>%��Y�2��+�U`��W���?�?�7\%� �7Ȅn�sʇ�"��~	�l����Qwʟ4V���yB���/t8-�u�m]}�%\h��������|�˟|�r ީ �\ml�����M?�A�����JO�%y&?�@��bDM�[o���9���Wq�K}���~ �#��G�����VV�h|�+��ZJa�G��8]~J�)lzՃR4.���d}���N�|ж�r��2����x����z����R7��<���N7A:	rhF�a��E9t��T��Η��'�뤴���<�ut&�N�WW`0>!3�wr�#����Ĉ���Ն���jiP�ldM^�xe�J��*����3	�
SpD�LC�I$NA�/����A�n��3�30(����.ת׷A�+��0}������m��Jˣ�_�q[)����_���g]�_0.o"'�tNy��-��(����Qk��o;6�5!��J��)g�J᭭m�w;2ڸQ>�r�Ƙ�����ǹ'�c~a�:C�+M��嗟��?�[���{�mqa�t�y��6Ͻb��!����̈́��kx�~Ц��?L�`� �;�󗾌L���[7c~y)N�>���јV���y8f.��Ş�x�=duW:�rG�������WO�!�y�q�ґ<��FH$_��Gn��X�ǚ-H]&7�]_b�oȑW7<�u�����t�N���:"��7E�jt�@�~�N�^������NWF������V;�l�Іp��cH�G{���U��Ż⎨����,�M��Si���_L���r�.q�S�6���!}�UP���
Pgd�G��Uq����O�I��1�r�_�&�Ԥ�&����'|��}�˲,� x 7 �y�k呯hq$
~�T< ��׹����t�o"�72B�@Tr��􀢝�fp5G�n��t�)�0���8<�N�K�#�`��Օ��}떕�U07�Rk��F���C�B⪃��?�m����S�i�lT�\)J����x;�5p��3�-�����r�#�
ț�W�[>�ZJ7���&#g��+�#׊D8mRo�Q�B�:$�L&�\	n;�$��~��3�l+O��@q�e�^-3Ѹ9�Y�ăW�)']�1�����Ϻ��Z�<�i��0�^�9�V<0�^�r�0�t�=zt�wL��Wm���_�E�������}����|�MGƚ�}�# ����-�&p�k��S�ۉmGL!<�d��G�ʔ~����6e���#<���{�>��*�7g��/c������O=n�{��S��dUF"��d��gBU��z�?U!��I�LP�3����#1�?uά���q�����kqB�ߌ�(�>:���1x�Ɓ�c�ȁ��-f1nX!�~+.ŭ�~�F�K�zC�LY��.ܔ;�;D!�y�z���t��iC�%#�l;�C��J�O��?��jJ�F{�GʒZ\����ɘ98����`{��8d�%���ؐ����Ϟ9�ƔȌȸ8��c˂�Boz�#2�˛%�U?�]ץ�Cm�~���K}�"��>���1���A����㷇�G��q�1�Q^Ed;���aګ�E9�ԧ⌃.Q��p@�5��]v�ɩ��[��4�V+ y��Ժ�H��/nd��&�O~J~Y&�v�!�;y����y��?P#�(>|����#���RA��#)oo�s6e)�B�0�S���.�Tr�(eB'�ߣ�����A⢄.O�b�L^<^1
a����{̱
�_D�O�s&�D���{��g��`N�4�&r�3U���C=J�A�t\GtXJ/�Lh���8��	��y�W�t��7[GD[Q���ĀOyơ
Y�z����@��$
=��]6?���a�͇¥��|�*��𠫲���SPz8��h���Q��ӏjP�Bk+���ǿ�����m?��i`r��Z�/�*2=;�y��J�G|�?�^5�s�q�L���l�E�K��=Q!�UZ~$;' &��yM�g�ą��ꕫ�P0� 9�d�������%ǭ����G��ͼ�	����v|��cr����P�B���5i�l�\�����pj���Z��{2.����阑l\��)��d��.a��?���$_�p�S��WZO?ڊ��n;�P�q�{��r��E�K&�I���~Q�s�8��2��CE�b��+M���y���9.>d�ΏM���Vl�nx�_��qlc����@Ĭ�oJ����y,9�1���,<�IVj���1w��4����!��A�]�s�?+A8xw�Stʸ��A�A�Yte�������8��n�x5�tI�� �m�$p]�뭢)�:���oB�#�+��Z �i*�z�o��WY?償>L~n���H���k�s�J��!��� ^�=(��~�F�����>�zj2?�K��4���b��-�����mJ��?
��F?y}G&��Y5³ ���d��os TZQ.�"�$� Z����
08����P��9c�*��`��*��-�I��#�1�*������9���`�%�wn<.`@���әIǯ���hb٫zeT��o��|+���H�-��IWڮ��e8�ꅍ�~@��@�ԇ�tp�u����+���,���J��Za�m���=��ӻ����>��a�o��>p�5�~)�/�'�&�i!��q��֖�>vByH�I!����gЏ���	o~i�����*cvfB�ւ�Oę3��ڋW��^��o��f���Kq��q�Բ�� �1��OV��|?��^'��p����c�<FJ�H]�?���0GV���7bT�Ϣ�M;�LF2U�#�w�E��J�\���ũ�Ř��!��Ʀ��ɐ��1݄��#񎄳�h�~;�^XB�����tȓ��տ�K�#������F ��1}._����N"gefOX�/)/΃��=v�{���Ɔdv<=17�2�;�;1�������;�}zyQ�ƣ�rxɩ�bJ<��BC�2i�EZ%��٣~Դ+��Z��{�*V[�V(�??
3�.آS7�.�r3SFq������7��J�%}�U�=�!���d��?x ~벮Y��<ʏ�.��V�[��<�범n�P\��ɍ��-۝|�e>�0ƞ�|��ԭx�> �Ǜ���ϽV�(��;���S��-�iEåe�a2�pA�i``Pq���~���p�r8˰��)r�IO|�?����v��7�n���/�痄�7�s�Б�a\$�G!�Л�Zǃ7�g�ē/�ꌏdh;�����J�>d��:3��0r���&�$�T�l�6�(���D�e����g>-]Pyщ�KUy0�%�t�*��J� �\��R��ɽ����5i6��xܳ�T�P�A L�P�2�����2$2�x���0ȇA�.&�-���_��DNON���H��A�ﵒ�0���X����-&BV�0��㲛�h[6�o�@#
|���"��=+WV�&�� �Q���#����8-#�ʕ���+/ŉ�q��f/����ɝ��gϸn~�
����6:5I�H��F��$%]ӄE_@V�2�i#1��U<V��X��V�i�*C�;1}p���&|s#%�����a�m��10�%�&�x��vK�%T�W|�%1�Yr�colSK������� -P\F�O54-�Hهd4����xrCu�܌�.���K�V�y4	���N����q<73���߈�����nG��rv;>O�А!?�vS��D�$�����u�뺊���c�	�>@�� W{�/+��!�7�3�*���+����S�<1�&0n"�Jz�c�-?�YN�q^I�ܴ���գ�=��_��4s\M�}p٭|�XFD˟�[�I]�W|�A �I���G@�龌m�q�+�}���A�/��zG�?g�Aa�&�o���w�����4�f簢�f�q�
�,��J��\����y�˯����a(��Mz�8��	��D ӦC8F@z������w`�N�����wy}�L�dz��M�%>yq�rN&�Q���u4���ԕ���x�����7=B�a�S�;n�E���L���e��"Ysj+�G�&��iL ����w�}C�Y���ȴ������+Ô@:u*OA�4����u0T�`�>!��|�,(Ɇu˚qM�H��h�>x�}�Y�>Y�������6J�n��<V^\�c�6`�1�bб�|Op���n^}T���x	1 �L^�JQU�Ƿa�ff�&cvv�oD���Ǐ|Lͣ�����[�9�++�b���Ǖ�N���I�;N���K2�(я�5Q�-M�"�^2�i{d�*z/��/�	��#�
F16x��Ge�Ә`��^�;ݘ�?�ɽ��_]���?#5Ƒ�K^ES!T�2��(��;n"�q3���������׋��������!ͺ�J��I�fa9	�M�Sy��q��f�qjb,Fe8�h�ꗿ�[�|�ϐ-/-����mU�H�vw7�f��̵k6Ė^����J�\Z�ჽغ?�w����H�'eTO�>G�|���8��+��7u��n�(��~Q�cNY2���6?���Q}�: :>����W��Q^�xD���
����r��g�2N��̇�U+�N�Q	�}P4��>&|�\ �u������}ol\�K+y�P1��8)�5ה�y1P�Vz��
�IR�0n`��

����O�?G�A<��r5E�P��知��]P�T.�xRI��{���O= �p�jhh�©��,�p�,G��H+���Dە?2�k��:5��S<�
(�;��A��'Zt|�\y�6�F��Yݩ��H� F�f���Z}�A��<S^�"��A�+�;��v�'@^��S��Z9�C:�A.Y������y�����M�����W��<#h*�	���+��^ ;��\W+?b1���o�js(�P*�y�NA���zt䯁��?ǹ�Qߖ���F&�T��+F+w�܍O>����+a�eP��$=����o��_�:��5�AC#�x�PZ�a�&l�@>Yn{ѷ�5ީ/���yԹ�����n���6�׽wmgwۛ�ܿ�d@>y�8������'�{�I�VX����CW��'e����@ʘ��ب�[u�6�����x�4�j�[��-�-�M�	�਌���f�x]��&��Ҽ:����BL�L{�bQ��0xR�T.H1��g�
��!�dy{c���R��?t�De���8^�ԛT�����d�M���G��'����_�㯾��uV�����IՑ=W�#��"�32�G4��Ͷ�N[Fl�KF�4�tc=ub9�/]@ n�1Y�>�uL���􃯪?m���~ĩYSV0y�/�Oz��4 R,��+�%�Z%v��/#���8c�.yË.�%�'W��'�cV�z�J���E�� "8�=�����r�v|�G�k�r�E�F2�A�����m 42?rJ��1�����H9�F���`���?o��2¸���;�՗_z�Y�Q�:�1B򊋼i�h.QG��4�'j��/��T��3(E��g���pSq���󪏮��� ��O�?T8�JN���N5n�h�2_�S����Ytp�S&y(����Y�&�WQ���<@�9�*WX}>��\�U��ol(�эF׻�gf�"��U7&?˟��)qH�B��.<�%>e(O�n��OU׼���:��8�rs��y�iY�8�*=��7e;���5�7�U�i�*������P���9iО�O<Y]t��`�<�/?�"��~�炍�����P��2U9LP_��tɃ��ۏ������??��gE
z���G�m�-���M�,>J���m}����PV3vw:���A��U��nW�Y'�d�=z�$��7\OdnGNJ���I��������?%_u`37G��(u;jF����<�p��鄌��ή��ɪ���b,�8!�C���e�I�d��E��������R?*,*��}�o�&���ͺ�7m������ʧ����b��/��o?����1����v�U���bL-,���q���F�������>������҉�p�d�I�2��n݊�'ʿ%9����B��t)��e���(����G�_� �B�&ɰ��
�.2��j���q�Qd(.۽�%y�i)Gd�yj�l�:�Z�3���-�J����tp���9��t��m�$��k�o�S�����E�'Ӳ��ҟ�*��K~%��G�eA@9 +j���Gq�̙��{��F��:��[�n���Ƒ�ݝ��qJSq��FYkK�)���G�I�_@0W�AW?�khI�]�#�����"�]�f�O�g4��M>���rف�g��Ғ��� _N yL�����EcʸC���|g�<&���fi�#GY\��gA-������.q.��+�l��K������D�?���L���L��A��-rz�̂N�t�4@~���A��G'�CX�2dO~C���q]�W��qՎ�k��_<����-0��p{+Y�%�p��������g�~���,-,Jjy׏�=&=��U��Ld~܀�����/����:�����d"�2��)�q>/�x5lb�{W0���1���}e{6�x�H���'#��ݏ}ՏoI��1���Fn{kG�؎[���^8��$Ϥ�����ա����RO�dX�����E١����d�*%������9;k�g`�ܥӧc��������%?��i��2��I�vǕ>d:�>�8����8⅓x�x|�}>�N�&��e�񋯢s�f���1%c��AY��:����R���?��{�V������/~���dG���{��W_���_�PgG�ڇqAr_>w..����Dm~<��Sދ74&�{\�A~�H.�4PW�?�7uh�?H���\��~V ��/��G?��Z�cY���~���q���<9~�U>��4�8>~M��(�Խ4q��U6~#����]�� \OI��2��+�d	���c��f��yd�R�9^?�'���	�1�r�'ߟ#� �0���6�߿ϊ�D�2[)���0����bYIR���Fi��R��#W�@]��B��9j�<�5�.��.=�D��W<O>�:��Wf^���3pV��6� e�q\+<�h@ #tZ:��+��i6|���XTt���p�������)�]}&TÅR�]�/�$�rB� 緵��"|��I;��Rw�2p�j����X�.#� �V�� �7�Jcr/?�e���b(��|���M���'w�q�k�p���2�O��ƚ�j��w�ɓ���ό3;=�wEӲ����m)������	*�<���EA?��QC��z;���������!A��@�ʧj0�|��j����]+�&��U����q_��E�7�Hg�+[�3�����ǒLn��zɖ3������Ut�t �7��L��Q�F�&v�/�����T,Ls���
�Q��ѣ����Q�xL.�ǐ��fJ���cFz����u��R�6�$LzM� a��
�qT�)����������'|>Etp�^޹ck��]]�a=�z̞:��.ǉK��hs%n��/��~�k�q�x,�V6���_����&}�EI߆԰|]\���dL--���\<x�$����xt�~�����x�
��D<F�#���j%<#���e �gT�|��x�M�s|�����1�I�!4(+i&�2��GHW@r��#���/�����lA+�΁�7ăO�ϑ�ρ�Y^�,������%�ڗ�UBF�.ԪG�������<�����q�P��Jq.�O� N��}��9B��s���zXgԈ����NKcʱ?���N*B|m��"�00��Y(��N'箓ٍӛ��Gb_1�$�b<��#FZ��8iڝ=>|�$����Ƃ2�<P0)x����
[8&ىT�����0=陚��%��]}`�ܱ:7��5�{�<�����~��]$Y�SGh��Ӗk ��Ф{D�(D�$�
7�	�V.DT��U=�����J��P3�h*���m�iY���Q"��I��xCo�7�ȕ҇4��3�8ɻ�� x�������&>U�#N�v�f|����N�y�^���U����[��wN���.�{����#�59=�圥�����Vyp�_�.�}Lj?�\�y����s��g?�����#��B��Hv{��'��������7��y���)���	�Q�d���?.�dB���0��j@5�׽\ǚ�Ǥw�P!I��Jx��	��N�mm��n'�d�u�wcgs˛�''��H��9P���G��2�X9cQd�ӑ�&�-o�����9�azDSz�07Gȕ7	���q$��x���ǹލ��)�� ����8V܍��'�9����x��t�ɞI���GƳ�����O{��.�-���(cP����G7��~�c�'5��iZ`��d�G����S~tc�|ȸ�����=؎-�wd�vU���l�N�ǅ�/ř�bD�҄��=��ڎ껫�k��y�v�ݿ�ƪ�^����n�(Ab��FVVc�׿��_�[t~��X��/��ǿ���w�B2��=�v�>+BⷃS@�����a�g����S��9~a0��i�p�W�1�L�1~��s��֣M��٫c�#��
5�2>hlT<� ���`x�1�L��C��;�#����U.�6�<��_�.<o�����[���~�J0x����N8�}�;������� ������5�N���`]S���j����Z��;���-5,56
�G�<�HAp4� 0�T<��2�ƍ�*�_�=����~��p*[2K|+��)�*m���Lt�����ɲ\
етn+��9� a�;6��g\���I>Gy� #��2�������tL�6T?�s�E��G�A#W^��vX�R��ѫ��%}�d'NT�'�0DJ�R.�`�78m4)E��L���	��d`�Xȁ�D��'Z
�:�OAr������2Yj�i�6�tt6M�Y����x��q���bX���]
~�!y)W��D ��o���I#��+��W�7��%�Na㐘2�5����{��I�E8~L�;���^"j�Ɓ�ePr���}]��L$��� C��۱��*џ���������D)��F��d4I�cgdS��S��5�*3nD!+/��M�h�c+���F�u�6������.���q'�9y��w�\(w_��M6R��a1د��P7d����0��:�	��ų2F��c(V4f-]�W�z+�O�r�����ft�cC�����Ա��g�9��4Ie#c(\qj8_�W��v'(>lH��� �d<�H��G��U�i��_Y��NO�/V:1oB77[��ݍ�p�f��H7)�s�15�ss�����ɝ������1��ݍ͈ݝ���#�1����%	ƅ!�qw7��܉G}O~���u3�o݈�/��#̡�]��P���)(���Vl�����Ic
z��!���/�td@ޚG8Î8�=�~�Lr�1���� �F=�6�g����q��J��Q�w�Or�?�Pn��n�B˜��.��G�R��q.�[�-�h?�ࣧʨ�h��В�gc)���oր|�c\I�H�F�OU�,p��:�帎d�_���k@_h�����x���j\ e-�*/�R@�J�`�N��������|¥d�SKl�[�8�+��-�We���R*�ݡ8�;PH�R�*����6�3!ll�0���d<J�|����=Y�U>ʑ<4 !���˵&#E~�t���6��:��a��ρd���X��.���I����e�3[/�;�`�D���&���d��i����;�51Ĕ��у���5(7cw��:��bP1�U��i?じ�(���7pۖ�J�<д+e;��q�D��$,��@�ݯ��I���xlG���'�^����Ѧ�0���F��K�qU�m��h���ϩ��u����j�:���#�ɕt?r.t��ᝫ�ir܏���w�rB_�	�ίx�τ�!ƞ3��|�6V�06X��ѯ���|4�����߼�7m�\�K�O�=.������'qLoOr���%�d=�2P�DwX����_Iw�4��Lp�V�#��H�#�x�+�f$��̛>���4��;�f�ⵣ�L0����t,�<��'Tv�B��g�toGƂ�|~Z�佹G2��%Wu=Ę�~𕄍�vt���v&s9�/_mon���j�>~�Wc�Ɲx���c���1���v�=(�6�.��ƍ1lL�bem�#���d1�+�	y%��i��L� y�Y޺R:�|�K��L��y<�F��iIi���*���8��x�W�k�7�+�}O��d��J/��-} :��%Na ~�G=rlO^������2i�q�R����M�U0��_��=a44�@crǽ����{�g2�s�/MB��/�~�� ����{B)��7�8+8{e�pO���2|�i���'~����U.Fa�U^�e'U� I�u�A$;i�c*�\[��{��T2�9�?Θ�-�1���vg�j��#܏(���ul��$��p�3E�	����D��+�@��ơrSo�6�LA2�	xi��gs<�2����q�9���1M�ݮ�G��q��bHiɞ��Oe�*�	��� ?Mg��(�d�{��<�`��YB�L�.A�890{0T�1i?�&<p18ث�ཻ�_~������C�$��#|��WN�s�;�(� VU(_��21Ѳׇ���*�NNN�����E�eI!d�M�sG|ĚF�S���x�N|,��Q#J�D:<J�n�m�%e�+ ȟC&��no�G�ʟ���cb�2�#6�@�>9�G���3Բ��c�Z�"�1�1p��1��w��0�a��N��s�cva.V>��*�q��%�y,������j�;A��n�
��y���t�ׯԏ�7Y�S?�kNtu��Q�vd��>��u�;<���a�af<�g��?�1����M���'��͍��Q��D������I�6VA���������:x��WeY�169�� �n�����)%��7�he��	�r��׊�ls���ɧ<�d�D�?��/Ǜ����Eȴ�3:�;�S�8d�����e;�J_�T^�de����N-�<.W�C��k�8�x�V�(�p�!�+^�GD�c����Ʋoql̯�U��A��O�?Gx��0��=�n޺��|g@�����RyZf��H���� �I�Z����C������b�_�3`�W%������Ɂ�����S�]���~�Ho2x
�/O8J�r�qJv���&mș����\�u5>��	ȈD8�(:��.ϓ�~��M00�Ln-�:�|+��g��!��$c�CY�h��٭� ��"c�:�G)�{L<�P.F��Z�j"Y�[���x����~�n�i�az��������*`'�/=��Q>���e� ��i���\q޻�(x�:Ƅ}a� -�@�4dj���a�D��&#Ekk������0=�Y_�ƀ�a���.�v1�����#�I<��+xd�q�*���T�=�����8��<��&cq$?�GepML�/��T#fd�Lql�&I�q��sZ?u����t�	��b�gEÐ�^�Ր!?�F���Cb9���R��+�\���	��5���=7C�a�kH��w���'��%H*�p/��f|�����/~�q�omře�~jB�����<�юj'8U����(̧}����g�d���N�';q�����x�	|3�����?�WY�2|����v�Al>^�M�︌�Nw[�%#�e�j�ѣغy;v�܋�Ç�Ê߸�vf2F%�3����+��tf��#�w�|�����=�;d(�[ҧ���|����!�?������ʜq��M�ڔ�B�c�R�]�8�ѻg=��A���Пw��ѝ�3/�a^H��^Tb�W�����V�t~����(= |t�g�)]p����ĕ+y ��iw�:���/\вo�cS�2-� FM��z;�r�q�ײ����7�<�Y'��2�vܿwϖ7��XQ��F*j��@��w8ѿ���t&M:�`<t�	��o0/�����Y��&���O� F%�I��̃��	��dgP��U'��2�}.��7%�ym�H*\�٣�dA��/GzQ�K��SF�2B�86��m����,�inO3��%�f�,.�`C,�59�M�a!��N��po�G����at���]��?�[��g���ױs�nl����Fu�&|蕌�/�N>�����T,�����5 ��x�A�G
3I�n>�kE�2��r]�����h~��A|s������RP�(�_>l��@�����vQFm4�.��	�+E�8�`��w#1����Lc`�ǚT����A��R~��;ɛ�~?���H���P&�sҀM�A~����|lΗ�$zL��X�\	tX������ʃ���(�Q1�0�X�����ti~��;6���G�oD�%����xx�f�>Y�tc�1"�ҟʸ�ͧ��Q?�lZ����j��9��+7�jz�� �|ԫV��_NE��	�����Dtddon�����mM���f�t��M��onEW���;~arrL�#���b�ĉ�z�jl�q����Q/���C1�'�>��Ǟ!�
����_�͏�N�6Dſ���.��;m��<g]�?"��Q��SGtR�+ɦF�ȳH���r���4���~�o�t���YF���Yp�����`����Eg�~ϯ���_�7��Q�&Ѻ�<O��>�����#~���g��6 o�.g �y��������XwWġ�\`�qC� SV�^ؔ@A�t?ï�_�_��0+Y��ҡ���ke �lđ�_�'����\�E��J���m0����Λ	�gGHH��I@�
�P�/�٧�q��E%e]�P���rГ[bU.��`n>��s�d�M��`�%d�V�Lb��IY�"M�%͆�~��$���x%��,G�8�2�����l���>���	O�v�V��W_�ڍ[ޗ2��eL��Knw�����W�l �LOK/G<�3h�ņCx ����mFtsU>!��~HO ��{�'��`!�hq������5��Ǧ?{��?�M���X^�=��th3��x�1|#�`fv&m����c�0�����JY��Mƒ��Ȗd�ц��炵�ٯE�y	�4V��T����a���%�����W&8M��`	����!��+�]�_���i��R��C��[�g�#�F�p]Ox9V����F�Lg/�ww,w�/��u�-�;+k1���ҥaS�O���|N�*w|b��Ǖ�����Ǭ�3S�������vU�2��C�.�u5B�o�B����Q�*�ߏeU�c����V��_Wu�O���֭;�y�~KΈ���4�q���ᮌ�m�t�k�N&�_����uWڮ�Ԫ�_�˯��.�������ҽ-@��Q�/��<�8˰�@?�K����#�a���]a�V���d��1���X��j�/�j��U���f��=�4�t��t�	餁Ky�qpi��׀t�F/�8�Q��.��(W���9�4ʹ���ƩS�,g��l|�1L��Aޟ7��	S#H�ȟ&x��~ܽ{�k@�Ђ^���˿�Q�x���Wy�0��Ap�~�����*����������[�1�x��%E���Z��l��goL"�A"�¤�[����r����5��̛몟P���!��z�_%��*'��dؕʁhlb�hD�R��L�6�Ւ�0���Z���">�R�x�s��x|G��X�gL����m�IH;��sq������'q��c�eDF"�ޮ�ⷼ�i�+<j�(a�K��C����k5�d/n��דɽ
�m���;��!\4�_a�E����3&-o^r�$?r� �'������]~T,y��mD[�-F>��##rH�(fK���wӘQM\��4���ŅXZZtY<�Aw�40|ؤ�0ڗ�4�"��C�nw9V�����W��Q=Ґ�H�6�_t	Ȉ�%�g��ŁUL�N����t��q��%�� [I�r�|�^�r��7 �1>�=���qt
}�UW>ͽ�q�����%�Q���I���$���0�� Jt�0>���o���w:��a��&�������'�늬������"&�9��/W׎�����IY���Owk7fG'cyr:��mu$59B���&MR�릆�Рo�ʏ��a��Cy�|Cu�p6���/��?�����]\���W�D�~3��?ԥ�F�m�N��M|�ܔc�1�j�͸~?�K�
�+]�d�K�����W�E��@�*�9۠W�oeWm��/���e��e����S�Ȳ��_��0��h��@h��<�L�Y#?�ꡥ�j��ĉ=:E����5 _���~ {�Ԉ~*ɱ0>��Ѓ5��o�j�TN�k)��i�Ci��$��@�n�VTy�l���YG���
��x��[d_�3o^I� ˠ���!��A��L2-��3�c�O���)��|�H��M�� (@׿��Wt��H޳�rT3م���$����2_V)'82�iv�,�H����x=�x�Q&�ñA���Xw�Н���Py��
g�(/�9�u��cP�Ԅ��	sws�b=�OpC�A����2�4�O�x��1�a2�+� <��+&+�?��=�:&���4q1H02ܫ��w�=GL��2͕���9��{w�z5�x�`౺7-#ӯ��Ǿ*VE0*8A?�5�jrs#P���Hf++2`%#&��a(1I����c���6)����&�	��%ZL.�"�w��±��Gc`쪭��#Lm�	o��;��_�Ϥ��~|�|��QUG��^Sd��0 &�A�JQ@����a(�+�x�Hm4����mB�0Ƅ�����f�����~lS��x�/�����8O^�R)SUS��.p��,޺���Hݠ��ӿ �d ��*ld>�yӰ�Za�a;M�?u�D,�X��ى5�dܕ1��îd��q^�K�b݁�b��C��TF<�6�'#�OZ��H�w�d�x���3��|>J�Tn� �T#m���ʨ>�@�s���iC�+=e�a�c�h9a8_�9�~%_ �g��s����Sz�t���HzA�M��q�c��A�J���C�F�l=�Z]�\��6P |��7b�G�-�ܕ���*�i~<U��U����=a�b��ǝ;�cc}��U�X1�U��N�Xt
gx@v"��@���x;��x����o�K��n��ge4/���7�)�I?��a�����S�At�T�K���e�ʓc�S+�e`�,���Tߝ̎���wxU/ʂ?�>UfV������V�\_az L^zP��#��$�$����/�t��hh�ۏW�$3�F�����_w�H>?���yU*�w�\9�A��övw}H%���&�o$֤��8ydHL�̊�&IM��/Y����XO������3ڔ�HK��s��Fi��凈�q�+�EubO���z���z���7e`���x�jl|4f5���Q�f���Ű�W��[E:GBlmm�6�O�	,�%���ظ¸����3[�y���H�:�~���1$�$>e]��7��J��\ u���_��a��@�0�8�?ƕN�Wph��X��ܗ�ñ2�N�M#2Xұ3�qf�D�틗V��G������q��˖2�Ƅ���Y��3�򍄳����H���I��v�>�1��P�LϺ��CX��=�$6{��}����Sq��1%=XS�jw76�;�����>9�Uu�������ɿ�(I��:=��}7N��NL^�Ó�2�gLy�g��'?��6�6a�/���QO�L�{��������R6)�4�Z��^4��F��.��1��]����R6~t�+8�x'A���2�����/�cϖ�~�QW½��[�P`�P���N�S��i�>�Jv��6NaG�{� �S�����O��s��O��N��}7��;�?*q㨱=�ѰB/e*p�)/X
���tQ�Z�v�� ��t+{�hy����ZY�X��#lPTo�uYܡ�y��@��i�1��D�qA>*�gA���-��?4����w���di�mb��ăJ�˵P������s�W?b���9ڀS�36=�.Ci����F�`��ܥLy,��Z�8�tc����>���/a	W2oL�>��I���D�iB|��kqI���^G���V�����٘?y:O����4B͛��-�mR.�{�g.y��q>����7\�����0@�a0N*��'�䀼H�w﮿�J����b�o��N�0�1 r�1��6�[���2�*��&h�X���1���q���B��N�"����]��1.��x��cÿߺT�rчz���J���m�c9���c&�v����2�#�̳%Qq�����NҖf(�{#�⬟�4�$`��j� �K�9aN���K�bh�{�1.�B����c���O�6��D������]�����������=:���3h�<��_�C��7ǘ�����8�⍷�y3��Z�Kn��t�.���3��xr�+Y�j{V���&�n��䦎%G�A�7�>�Ϲh��#*,���ob:�^��{O�1v�n����,�bs�+�w�t��*��(^���e�P��
�~�2���ү�On�4]��X��~8��y� ������C�Q4x���*Z����U@��<ac>�UK'˧>�롰�$ɮ�G��S�� �t��AV���S0�W�}߼n�x�����~##lkk�v)Z������j��26��P>�
� ���kY���qu�Q(E��M�[Zuf@�yUz�=Ã�T�`ӑ-Bʓ.�Ȯ������P�e1��&2���g�L�YuKِn���G��JrY��4H2����.dc9��<�i�8xd���Y�_�JA��7nƗ��(�=�q�����9>��P��}P�'N��s��쥋�|rɛ�ǅ��X�#M6�넌�aݥO.,i�4�G:��d�$��B�Y����� ��M�4�w��=��t���(c�Rq�;�;q��M��y���F��/�%�m�g�N+eЙ����)�|0���1�X���޴���6��N����TV����$G���_����� CfH�Ǔ�#G�,�>�\F4�AO>*�չ��;�F%�c� �|Ԓr�L�7;���\�iR_T�^V�|t�]�qp؍��mű�h�@��� Y�W�����	�O9�8>.��J���?�0<�O>GMu��x�l�f��L4��v��~?DWӮ�3@��C�#�G����_⅍�{J�e���h��_��|.^��x��byv.�҉}�#��?�	]1Zyĺ3t���֡ѡQ�#_,�M�jǙ�x����w߉!x�2H�G��$��=��n<Y�5���sB}�����d� 6����o���8��䋸�Ւ+�H��Tz����2-�O7�'�?�=�
@��"}zi�je���9�h��l<�?xr�+�04x��q�QAh�E�a�M�2���?�@)��=^���'O��@��|�Sf��<BJ�9����,�Fe0DYk��B6���[~�+������s�8�+�YƣE��(:h`)
�ţ������`U�hq$�l�P��;�����p�hq�/��D�:�z��_�w���X3/a�:��U����-p��C���t�NIi2��ha��껥Q��rɛ�
ɋS<e�8���~oeAh8���7�X]v�5���f�^��)���+�ժ�P��|,����b������zl���ؓA�y�Vv�T>�w�jbք��߉�鱈��ؙ��p�\,�z-ba*F�9�A%u�b���ؼ;�UL��丸���7ÆG�bltB����L�n�r���x��z�Q��۲�5�4��4V��6[�a�M���P3x �D��ף=��xC���0R�������#2\f��n	�p,{��eadq+)��a��4K��1�	yzbTu�����e����R7�7��#Y�i2�������H�h�U��<�\�!+Q�I�r1,�e�}�狱��� �
�+���7	���ۄR����4��U�W�`O��5��r��|ل���s�P��+|�2	a���p��*C����E�|ΉzKicB��E���z�����f�yy�s�#U��ƞ�ngo7y�7?��x)μ�jL�9i������������J:3J���UR2�$.C�FӿW����U�)�:�v?�6��<Hr_6�ڸp��#"��臬�avއ�=9�.Đnf��o{�7�r����{2�Jf�ex�����X̟9����QOPza��`�}�lt^�GO���TL��3�2v�WW~��q�����?������_������6�5�%��c���0\�_ҠɱG8O�.�;F~�LP0?��߄ER'R�5��&=�-}���=e�x�c�tJ����|����_L�ޠ]�A>mL�J�f��8h7�p�\���8�Ե���p����
r�)Ƥ\���A��]>�<�tp�ck������g��9BJ�9�#�D��&{:��H�^c=�^ՀP���k�A��jd���1�t�I���sO\9p�O�St��6��'�6Ȥ�t��Gg�+_/��M���x�׮�W�����8�nëM��]I;p��&Mpp�tjp�|�D\��z�:TW�3�<�{���3Sw�LY�5|��r��Z";M`�WQ6@2g�׼��ڲ���ɰ{�N��.zzc;~�yܕ������Ӛ�4��h����/��/�嗱�;n���T�gX��WM���ƫ�[�d5�v�Ǳ&�1IrZ3��e�
��a�g�9o�N�k�C����2����x�V|N 鐇��&��SxDv~�@�L��D�#�����G��Q��Q!{0��!�L�L0��0�`c�G�*���b���C�l� ���;4�S�ߺT�pՔE�X����l,,/�H���
ݽ���#C�8�/�0V�x�	�8��1)���oW*�����]2C�%�8#%� y��R���)F�C��*:�sV�_����߼��F��}���؁ܞ��>&e�����F��UJ2?�(����+Wc��i.��t����ȧ~�ǾeH_�Wqb>a8y�ĬN��V��
���9t�~/ ���T��?�;�HOcCaHf'���7w�G�~�}���lJ���t�8ޖ\6ucr8;^�o����w���7Ɔ���^�+�'_��
��k�1��;�~��o���"��?ţ���SY�u�׿��������oY�-U&:W���z��N�}��i����sc����Ce����_�c��rl���}��;y-o��>>r�4n$鯰[�ҧ�V�Jdެ��^��h<�n8�
���B�р.�Dyi���$��#�H8���ڋ2r%�"���c�]i�+<��Q@�h@&�[7oJ�9P�;զl(3�nd�������ACa����)[!Lk�n�#���r���=��2�/)qW��� ܸ�;��K���!��3��|���x�'���)y��9'(ǃ��eC@If�2�G:(ԽɜX&dc�-����2�L\�3)ȏx����쎗��>2Ȼ4����"G4p��#'�*@����o���x������ؾ{/f���`8:5ÒO�M��ذ�u�?�ً����ǟ����q���6��6o݊�[��hc+��vE^�q!�d���܌��]�n$;���/�^��{5&O`������ӣ�����^� �d�֟ gO���Zlnl�h����yŋoN8����AV<�>L#A;��WtY�}��D������#]&*mRx����d�?w>�]8�0t0L�9h��~��T�S���I� ���sL���,�2t����0ڠ�o�y�|ʟz�c+hh#��6��r˩}�<?A�3�v�cB�ה�>)ce��8�sH��S�|@}hX���=>N��N�|��:�2�T?��b��g��>s�A%'R��~�� �-W�,�)���?� �i���{"�p�YvM��e#2��>�u���=z���$�q���Q���M�[�o}�{����^��`�Ff��R���?U�{�$�~om#�o܍������/>���~G����f=Z��P��B�S�w�'chz�G_���K�`dW�67ԉz���7u��o��I ��o^��!�1���ق^ʞ�H^(0���Tc< n�絡�o7����\�k7����	�8�I���t��WcH�~ڼ����u���33s��U��y.�9"�~��ߘ/(a)�֭�+�W��Wbru(��w���#�)��'h�3]�<8������l �x�������]`�n�.R��T� �Q?��m�0����d#\J
O�x�	�^]3�,����y���&���%���`'r���Iq\��`�0�h�*��ym8f�?�Y�c@�aF��OH>��e�%�u�Jv����Ny��2�����M�Cq��vO��ĩS2���cg}#n��Ӹ�����'����������G�c���غ�07wⰳ�2|p���S'�����+��,(��x�MY�8�,teH�F�Ӧ�M�%�
��u�2,��ȏ�*�t��{�[r�}aO�<�q2*�GF$���;+��ڊ�$���<��(�JV1�0�d`lln�dt&.6�����v���+���Ǚ3���%8�1ɛ�s�'>i�+f\|x�> ����O_)�m�f�h2�'ꃣ���U&)�N�þ܀��%SRՇM��rT����<�@^�����cr� &e��D1�z(6ysp�G��ڃ���W�/��8�����K����3��M����WL1�v�O�*^�B��*��"�%����>�>�?���o�5�:�N-�ܲMC���Ξ>�c��x�����ݓ1y�{|y!~�W?���y+v��qCՓ���h�q��x�/>��67;�oߎ��������#�Q���յ�ڱ�7����y��q��<܋a��i>��>'Q�A]���"������ �\u�GӹR6��-��cI�79�#�t���4��3�7�}�%>��<m�L���wT���?��G*��P��j�.����8�)�|PG�U� �2��1ֹ��:17;�����S��,|[<<��#� ���Y�v��������K��6d@�� +�'[�?3 ┕�������lԁ���5��A`�NH�
=��1�?��G@<�3�Wp�i�ݝ��x >�̣ ���<�k����G�:�@>:_֕���up�y�o]�.S�-�ǝůy�B =�M^̫�"<���ܥI���A/y�ŏ{4Is��YyE��`/��c���8Н��Ɔ�f�S�1��'_z)�Ν���y?N��X���ףs�^L��đ��#��߽�vu�>�	V���UlL����c�G����U:��D/�|������A�کd`y=�ӫ�K���s������I�=�c�𱹞����ʖW4i�̕�q��@��5	�.�#�2R��glаY��r�oskSġW�8$�6���F^{��E;	aر:����4	��pV�F��]�{8��0¼OM|���#�|�LJW�'��L̄"�x���]e8����~)�_�u��NmfcG�}E��"��q��S���4��K�6b'ħ�Bv�:������]�1�,=<��79��%�����<~�d�f���3���`>�?t�F"}Te�x�"u�\qd�| �����?�sl��韤S��'T�yk��Ɋ�m��U�|��7�ÿ�˸���T?�䷿��on���ntv;�&��Dڛ�՗_ƿ���/��ױ}C7L�ᙖ&�������oLe�S�C���!~b:N�>��MN��C�$W�ԃz	\o���@n�y	$��B��&�� �~QF���"M�ks���+.�f�q�L����0�n?�r�o9��Syp�f�#i�/��qp�.[���mi�9���A��o��/z�>�������x~��;�mO����vܺuS����q)#+�, �qC�+�p�P��m"�'������8��N����h�<g�C0%�C�~��ݼ7�����������	�8�� ��L§��Z��Q/�~��M /Ձ�_�τ`	�A��%W��˸�����V*~�S�/�/�x���fd�r �7Wtxʗ�n+�x��p�u'~��[w����Ǳ����Ù�X��p������+�7$َǼ&�����{� �OŐ�8��x��1L=U�r������^_Ӥ�{�[yھ�`^���&^�h+1Ɂ��ǩW��Bn��A�@�����GO��<I���*�8���&��b`b��V^���&̡��j��$�t�0�����g�q���0�i"ƈC�x��3�Xc5��`�a���G��t�r��8��0�4i3���6��v��O�h���~�#�7���r���So�z�#�؏MGG�1;j�:��e���Z{��L�讜h�h4ɒ>���'���d�@>g�EW4�Gb��r,,c�b���lߧ���B���{q��wb��)���N76o݈կ��;�~7>���>}�d<�J��	]P_b���T�R�˙Ӭ��"!����R�2*#���Il�4��A��,ӕ���V[\}����o~�^y1��������7��peC����Ac�!��zp�vl>x�GObtc+f%�)������b�J��Cy�[�#�g]��{;j﹥�q�ҕ�f-Ѽ�w�U�T�$Sd�Q�<�e��	^:�A෍��S����	de�!��M�I�O��z+��7?�Vz��uV~�*�f]�C��w ?��*�zW��د2�]�\�.Z�F�����2��3�S_\\\j7mI���6x6�0<��y���q�ۄ�cX�v<��Jꕰ�PV6�h�Z��_�������U?V��m��H�R�U� �`̵�*���$@�v\���� ?(���;X�博rd7�t~��F�z�t9��NG�
R�1Z���������Ff�㢚j��^
�x����P��o�]�r���J�RtY5rJ�F��N��`�2�&�I�T<m!��oo��B_�x%���[��ǶVb�kҟ;s&�^��ˋ���u�(���8���|xk����gST6��e<q���97�ۍÍ��]Y��v]�� �t�TL��ƾ�t5�c��&�ؐ����e��D9n����&a��@�����O�����ܟ%���-��m���x���s[�B�,1�x�@>��*�X����M� r/�xy���cb�Ξs�E���0�`�-�y������q��	3�9C�澼��ǝ���Iv�rx�#H1%���e_�t��@����f���C_�� ��V�Hg���4�����G� �i"T9���$nl�s>Ǘ�6#^�ϟ�KW.����n ��#�:�43���{?�˸|�Z�sxm#�d�<������zt��(�}3Vt3z��S����P��I�XE�?I�g�L��Y]�[*�?e¨p�g���@�V���J]����JN�4���"��x���8q�r���w���_V�؉O��_��_��Q;b���Y��\]��G�cge5F%?>�4����9{moT�I�Ԑ�A����C�rW��=��#�f���oF��t��/���٠��ld��&���Ne���|�#���WЀV�L�%�,/u�����<h�y���|��(��`:�]����ѭ����&��Vt�A9\)�����w�ĳ�V}p��Q22�����8���z���@�g��p�|o�#� G(�{�ݻ����)k)�'Z]�A��!ݘ�U�����q|�JG)�����
�W~�4� ����3,�$c������t^���7;[�'�хG.�9IC�}��HcY��f:2TZ�6WŹ<���2p�����?��h�p��%��d9� q�/ڇ4�i�g%ɥ(�;k����A �p̀�tY�&~�v�7���Հ���;���f�+�)�d��o���9�4%<��x|���}�ī�㷠TGVk��L�AW�0� ���.o_I2�d ����t��B�,��W�8tr�0�/��L9��!�HO�W��f6�Rq��W�	+5����vwcU�
F�ΠA9�A��#�Oō�_9����Zn�R�/�8S�8o�(�;w��I ?؝:�[���1��˗���_�9	kg�oR��0d�lG~�1�)���e<��/�h�"V�yi�U>벐�f�l�19�����M`������Ȇ|�G� ��	§y�4G�{0'R�˗.ƻ?~O�}�?�,��w2��x�|�j������ń�y�V<������_�˿Ė����Gr�Ci�+g�Q���S1����G����^��2a���Z	�#���k��#���epS���1.Wt�q
`(��R5�\GgeП=3�������������}[2x�Y���9^d�H�%��	ڌ4�1��z?��=�iƛ=�7r�t\�˟�՟�$�ϝ���9.я��K�"�L��%�'����A������!��fտ�"�����5$�A�$��3�����[)Dx�Օ2q�V�I<QD�6�\��߆W��o��9^m����*�,�$�eR����0��0�4�6��O�`|�]�=���2�:6���:0i�r��Fc�MPN�[C�����n� A�v0^z~�*+ ���4p�؈��@^�U�N�ps��,V|�3(L��T��cb3�D|OQ��OώC\�A��AZ���w�O�C��leO�x�O��	T�=H(�A�Rm,�J-�����7��쁄�Ǡ �o����w-��1�4]��f�լ�����ގM�m���p}3墑�ի!�M��a�'+�}�^|���&����܈��?���/\�Jў_��z���~1p�c27���267��˱'��I(�䎾{�'��o˞�����뵗`0�8ڇ� *�vGެ��$�{�3��.\8S�(��^j`����G,��+�(yT�g�0r|\���8�r91}}=�޽k?@���x�c���^�ǫy�
c�Vd^О�^ɸ��xDF���dꚌ
& ���˳g��Ѓ�[�nIC^�CF��a�Y��ʪ��(��p�;�7."��Zy�=���[Ϝ�w����T�����z���������+�g/\�U�*��֯~k_�P�� Fw�c��@���_G%�q�Lb�L�����	=�����T�n�����O��_ྖ��M�����[�o���7�-��瘂a���d!�O��:��7�Ǔףs�^��]��8��!���n����.:sӳ�$`_+}��J�Q;*����HQ��U����q��?���71�ؗ�Y	O�����u��>���R���� ��1����)�%���g|�'�ۧ�F�o`I!���mTsiU& ?O- �^֭�6����T�S8iO�(����d�l�<�����h>���M�����o%��Z'��Fr��/sT��; ��kr+�t�~!���	Ho�����p���~S%�ꔢ�<Uv��o��pqG��[)�gn��C����d�ɦ:p�ah�HK���kɂ�WyY�B��Lf?eXe�vҡX�)BO���j�t�@���|��ey��ܥ�^��5�/I&������X��{u��$%9+��m�c����Ė�N<��qv��ݕ��z� ��܍����xk'�eA��L��n4�s��=/�-=F"׵�~�v�`�1��M8��U���HL./ƑVǔCy%MH֝g���upծ����R�)���G�ځb�˞D/�L޵յ8u���+�}��.�ж�J&�8� j�%��uc����Cjnn�uۖ�)cj���i��Gf<��V�Μ=�S>����32��8YҟU��I�@��oȑ_E̫Y|�����2����/�3���_Ď�>ʡ�%��a�!xg�F�I����F�$�[�Nʺ`�H��66���S��{o��W/�
/|�Mm�h�J_�#v�t�:w�ǟ|����Wr;������SG�{�ow�ݍI�w�h8:2B6vvbK�N�>/C2�����+��O��L��Q8t]����;�x�j&����Q��s������lFd(q����4��A'��:�|���}pߏ��$�]΄�h�)�����S2N_뭸p���|�`��n(K܍I#��-������_�E�(ρtc�#����Of�����X�>�%t�m)��_�)9渖��@�"P}�8�Hh�xs\���S�x��7���7�che�X���f���xڮ���׵�i Q}j^p�p
𼣟s~�ҩU45u�>}�0�I&��8��4c�Yi[6�ޕv�[��~�ʆs���8�`�L8:
���t�"����>-En�|���A4 Ԧ@.CeA�8B�R�ŀӣ�x g��3й���a9��'�S����i4$O �ϼQG��)[�(���^y�5���*��^��K��8a��DM��F�'��g� �$��K.7c��1lK�qЈ0V[�Dw��ƛk�G9�ྺ���FT������J�m���X��!�2�Ty���<��vv�-�m>����O��,�&W�XQd���š���]&8�T������J����r ����Y�4zq�`~�q��L��VFGU����K���V󈄕��9>�<eZ���a��/�-�.^����`|�̙�r�J,�/��[7�w��1'yB�v�c�ڽ��L��>�F���9�xa�.���S��y��rtx�zq�*�Ǭ�����jܸy���q��I~2z�@��4n8AMXșr�)٪��V嘜�+9NI���o�]���+q�����_~Wb�s���"b�X[���wcS�,C��8�)O��P�
�ࠠ! �{�ʸ��N�Ȑٛ��1�c�f|���I\)���x��:d] W�l��j��Y�H�� ���MMr���8̉��1Ë.��20��ƽ{�Q�0,���Ԅ���%�W.����Ǭ�2��ܹ�>�U����4��ucwq2��3.��_���o���+q(9t��x�o�W�eT��ڮ�9���ۦn��W�z8��@� dW�9rl+���cz�'n�єc� y�����־��쎗���H��|n�o�i;%ׂF���
�����C��Q�͙w�@�r��չ���`�	���'����1�moo��;�����sïZ��*��F#-'�P�,��4�i��Q0��k�V�B�P�Aŀ��C�p*_�AT�]���ޚw������ze�
�	g����9 �}�p��,
����W+ׇk��/<%/i^�$=�)�#Mh�D�j(��U4o¢�U� ������� 7%%�"n0U���g���Q&Y)W&�pt����F����$ƾ�����޻k�m�2yKp�ǚ�9�GJ<��g`tW=��PD�����5҄���Z���A�ǎ����yT�{�>����kW���o�$ϧ�4	�6�u1�w�͠��mB�D��ו8�|�����K@��Q7"��y�>�+Q�:3�` ��q�5d��'�}��X	˽]�0�#)Xq"ߔ����G��;{�l\����
��d=�ly��	�ǆ�ZYY�U��?vܒ�0E���B����-�-#�o��K�Y�MG&�����Hwnxޔq�������y!�U���E��/}�GZ�/D���N��v.�i;G*������~��ވ�������1��S2|V�ĪodnlƐʟnm�#(�e\����G�U/iaL�N�(��M�(͎�1&�p�<��o'J����HFs��>���۸�:d� �>�K��	��OC
�a��~�E�hl��D�P�2�X�W��CGqbf*�v������ή�-}�Z^�s��o��G�«���;2J�ʭ��{EyOFؘ��Ѿn�T.�ȥq�o~'�~,��~�^���I���YɊ�zu*W���-qەN����>�x)#��O�G��g��G���^��4�~�O����O�\d�@�� ��/5VR�����A�y�7P� �4�4�l��!]D��2n��S<"&/uוQ�s�3k��Ve�)p�T]K��+����]�7n|��4*���P5и��k�A��(Z�9��R匘�R��W����\�\*z���倕f�dy8�t����l�J��ή��A7m����O�pytb��<��C~T����AxP�s���ԟZ!Vv�����ch$�JS:��r�77������wkp��ߨ3i�Y�rȜ:28B#kH���9��f�=��C?�j)˙Y���Ky�+`L���a�!4�8����NLv�bB�>>���=M��� ʢ���at�xlr���7�ې��'�Ӡ�#�#���~�ّ�'iӄ����/ž��w��p�8�@�0�I�o�L>Ց7 ��?�Q��9��ȃZ��iLe�Ys�\%�^	�,�B�ohxi�p�ߨ;��j���^ތϾ)>{4+å���=OK3S�>�O���HZ�������r����X<q2F�e����R^�r5����o���6׷��zT<IOx�6-���'��㕸~�����O��kC�Ԋ��k&#lG����ނ��2�\t��&S�H�� >��ۓ��rJ�o��	+P�c��8D|B�rF�D����T�{�^y�j����O�]߈�������>XTd�]áQ��t��#�o�����M�GF�g����ڞ�VG�2fdd��c���r�{��8��{q��cD}���#���}�:0�4V]l�Q�����kd �N����A�re-�A�������Ӱ�HLȠ�$���461���x�щ�����������q\��g_~%6�lģ_};_ߋ��V�v�U�#j�����^̾�J����s\���W^�ñ�b�:�|e䨾�?9��i��y�1��dY���#PcS���6�2�+�<�-o�!
�>}^i�T��)�Sr���FSk�'��ڒҐ��U�yn��(��O�9ƶ>�4���^�a�j0G՘��"4�M�6����|G����zϰ�>QV��K���w8._rO�����A�.R>��
T�{��a���{�1����e�G��P"(���p�_�8(�P$�qP8��C�,�]���J��ah�������v�
���>����f���_^8:����?qJwG�u���-%TG�[P���]8����4p�Wd`�(N��0`� R����Yw6{s��4�_��!���`�����&4�Q�Cv�+��A���yV�� sEUKe�ĝ�� Eû���c�����]M�w��o?����(V��*���w�#�1�~�#hM�|�\�ɑ�f#/;��4IhU��'��r��L�0b�_G��������p~��?.v5�b�qlư��G��x>d���&�QcacIFѰ��n��84n����`�q[� ��1h	X-Af'�q��q{�VWW�F�믿�s�2<�d;�� Vyī�eW��8c���q�o1*c����1V
�)�2)?����������_Ǿ�Ǐ�g�G/ Н]��ېl�f?mO^6���W�	}\[_��Dt�:��=]ԏ�&S& �B���~��r���Ab�LN�'.G�&2e���9�>EX���Ϋ���ӟ�O�z'��^���/b���W��M`LK���G�#|>,>�6����������.1�Zjl��w,�vd�;�{+^�ч1q���	���v�x��P�Jh�(	�ץ��؀ ��f\�3�.x��~�Ƶ1�	YbԠ��*��ℌ�c�7?�TF�a��|6�\<k;�q����ǿ�$:��:���<�m>��J;���X��_�w�ӿ��?�QHG:*���M�d�H;�4F�u�?V(�jK:P}��^�9������G^ ?�~�Cq��2Fd�d�J�"�X�D奬4�gS�&�i��ťԓ'�s���l�f\e~��(`���,�|sX|��V/�C��lW��*��B�ަ#Y�e�#pK�����U�)��O�ϻ�ܯ��܈�F�ɭ�7�0��y)��iW.�9>�Ã�3�8^4P&�[���2��M�+�P��K�k&�����k^��a
̇� �����Z��OO^�I�e�4ش]������p2�]�|�O�kuL��(�	��LLV:9ȵ���뤼�9�����2�L�T�Eg�e�#N���rӏ87��0a9�d`q�<q"9>�d8��K��{��4�l����qL��]�&O��c4��q�S�>��<�L�8��1��c��b��W₌���g�#91�k �� 6)u��W�d��Ǟdv ��T���H5x�-��u,�����l�oʀϋ�.J|�|����Q����/���1�A�����K�%�0^�%:����(	&���'?�N� ���/�_~��7����*2!l @��(d��G��2>~d#c�O!qe�o\�8qKq�JQ�V�Cs�����7A�щ�&�U& �gY؟���O��'d�v�WRΉ^�����p�t���+1+���W�cSu�a;#ꘉO�QM���bH�1��3�s~�8=6����q���O:�}�<�����嘼v9.������{���e*ُ8������v�}�@Ӌ��:] ��\W����f>����P�)�*C��]{�Ҡ�X�tn�pSҗ��Ŭ����L�?�_��/����x���1����u,#��suC%k�Nl���y�����ę7^���d�O�K��$[��8c����m9�O��n7��T�1�x�m�¿��W���(y#�^�V�g��e&������K�QH.�2�\�.��/�|b�������݇�ʏf�7u��,/�/^��cHS�������d\��|�GI���Sտu��T^����4<������ ?�Ǒ��tv���[���C�ꚓI*Q)U)y�oAw0���P���-| z���3o���$�%��:��_��|����A�
��d)��?I�ƶ艦zI򞜁G'sy�L��ɇ�$6:tN�;�'��H	]�&~��*�eyp��`�wYY6eV�է~�+����(��6�)��	?Y��RT�m�j�aO�Sb�>?�Piq���xF��|,�9/\����8҄��+�kOֱW%T�?��]�!�'d�i2��=1��I�������'b�������KWcw����)#Fw�1̛�ݽ8֍ƎJ��]��.�!V��ρ?u�o��� Z���� �:�O���0`cx�rY�;����]��L%�&�H��Yi�pW�{�rx����ɔ?F�� �I�H�h!��7�x�o>oln8�ǚ]B^R]ɿ{ �K8���U;�G�9q���#sEPY����/�7	�U7t�������ܹSg����F>���ĕ�c��[�>�t������B�.������Q���V��È�u呁/�;���*ߑ�u�ŗ�����%&�:�[��{ԉ�Ζ�1��`��s�T,��F\��_��w߉1���4�5���nj��/���(<�OU\~~9v\_n�h������ꊬ�m�tJ���+뢡��mHfu�~I�=P�Zw'޻�~��x��_��'_�\g/��yx���e��Vwv:����x���_b��Wc{b4vx4<9�ǜ^�V��8|�692I�Ю9��.��Թ�� X'��Tm��iԽn�KW��~.P\�?��W��,�'yB4�T�2��	�,3�C��1�Z=��\���Z���J��J\�?I?�į�w�~�Sג�k�t�7� �cvv._�i4�3x}�M�Z�>������Aww�oG�d����4��e__��@�(Ru�jh\:�JG�ͦ(,�X��
����%�Q �my�TD�U��T��8��Ƌ���h$�O�I��o�(�wO�+<p<�H����5`��,�ã��4yR mĄ]U����G~� 0R��;6���D��SӔ?���ᵮ�%��)?�J6���|��g�a�jء�x[qvv1gbZ�z����ǝ�,��1$�t�-��k�����Ź��$�;���|���X|�j\x��Xz�J��ȣ�'�b�3�6�c��ݸ��'q��bcw��j1x1y��^�Ӕ�Kg���TW8վ�*H9���5����m�Ǎ�<⣿]8Ο\��aB]�t)���]�_||�hiy���4���̕6V�0�r���&�&���짮�77oHG�l0���U0VTxB�W�t�o��������mM�j�Z��O�2qy����ɧ��F�#�Y��7�i9�.xư �K:r�I��}�
��9N��^��tZ�v<x� ���w�2��&'bF�<�ҵX�t1οp�+X+�������u�@������hc��?�I��ɇ2�_���%��%iRV,�1V<'��.���d�r�]��K�2���/q�^��<���G\����u���]�Ø���ʣ������"&�vb-ꎌ��@G���_�4����SL\�]nTx�E���y���3�<��O�(�~�E�G��!��Q��
�^��+����#o�)jΘ�234�A�|�A����q�$0�Un�D�䁕^�NgA�Џ�˘�'���7��7~��e�IFI�x��Yu�thP��Kܬ;FW��k�-�c5l�,g��'�ӽ�~0���u;q��/u�Q��� ,c���W�(�A������	���:M)	΃��+)���5i���L8���\���ʬ8�ʄ�Sx�ѯǷ��pN@��S iSo�R:Eu�d1&�3|��E<�M]��;�LD e�-0�a��m:��2|3p�PSzN^)O��9w�*[�a(�*�	�Nn�n@|�A\s�?8�'j���J��Y��U҈��E�� �x��1��ߕᵶ�oގwn���xR��՘<�,�>��'c���X8�o��Wicc+�����l�]�W?|7.��j��M���M�k[�������z���w���?��ζW�$�X��83g��{A�m��H�3k��8^���n��� �!���H���q� ~�r�[[������������ Y)�؉M��}�y\������t�K~q.K@��$�d'~��/�y��w�n���q�C��΅�AƤ���a�kss�^��(�d�+f| ]� Z�����d��ɧ��q%�jr��G��M�y�̅}��fE��AOK���F\����/_�F�[wn������⽿�y|�7�^y9���y����v67X�P�i�I0���ƹ�ގ��'�x-�TV�clRƹ�U��$�Pe��d�c�:Dʑ�<� ��ZM���]�i-������P���^��R����o,J�86���L,�?�#\وq�骷u�GcS���W⭿��x�o�6�%ߘ����r�t�6c��17�è��r�1�r�@�#�ny����{��U ԩ7^9&��ؑ�#o&��@&5g �ŕ��.�U8�Ad��OS a\a)_r��ָ�+[nSA]�i5�Py\Fx��?=^�L�X�Zu <�yTNp���N����	�\T��A� <UF�����7�  �����H� m�;��7l6�D�"�waN2X���T��P^Ҫl�� ���`~�������t�*��ER����a#��	B}�S��wELX�%byrx?��pI�*W��s�qg��f ��J�_���|�L(��+B���O޹� �D���u`� 4��.�G�9`P�9����8_�A�)�A�[�*��e ��\7�E�����C����_~��߉ݩ��_@;�!���0�	���ʋ�|��m��œ�To�V���sq��w�̵K1>�;����}�0:7�ƽ�u<��wq�����[�aR��������)z���������^�[q����8��qš;�W]M�t���e/C[r��s6�>}:._���26&�:�<u*� 7GD���n���������7���P@oV��_��_�~��[����nǦA&x-#������ʅ�`H��֭-�cE�q?>F�˷v�xТ/�˩��I����7��^K�`]�㘕1z�W��^�٥E����xL�b���W��%h?��!���rlnn�?��?čO?�Σ��y�8&E�PF#��ճd�����sq��~�1q�b��<�r����h��*Ѻ�c ���
��rΫ�S)ˑ1��%���􁆫hˣ�uH2NZ��5]c�!L��GV�\���%4:s�cl��K�d<Ǥ�������>�U�[Gtv&'bᕗ�ſ����W?���'cWF�:�Ψ �H�Re�#x4��?�|B�kx�R�'�-��:�+2�b̢�!�H9V���]�����,��R^�ϩ�M^�P���7��Ax6��e쬶�:��o,p�4�Ƕ0Vӧ����ո�@#�g*��\�CݬY�T&�֣y�#w��)�`<���ף�=��9�cOXzm]߹sˍN�S��J��PP�,��VA���gO�2��1���`Ty�isP,#� ?4��x�P�N��N�e$]�GX��W,I��Q*X	O���ա��t�D�||OB����/�h�1��L
��m�vRЫ��Ȃ�baq��5�K�{.����t��#=y1W����='@�����J����_��@΀>�	T��&*��a�{��'��.��j������]��7�$͞����l��j��rQ7�q�o�����x�ٗ�����<z#����%��=�hh[w���xSofn!���bGF���=��A��Uޠ�������G��=&H��X�6LBr֕�k]8���{��^��p�mD*:�q
����޽�O��Dnʧ�������W����x�7�W_5O�ja a`u�]�nr�?�C����Y_���?�oj�*Cq�|���Fx̛OO����rrC��km�mK<w�B���+�xr9&d���p���������t�l�>w>�cM��o������E��Ø�$xg����m����+����{��������G�t��&�4x�:�v�i�/� ���*�D�Ǌ��Y�a�m��΋>XN� �A��gpq-4p��9ư�D�@YJ�l�5r�^q�c�	����x��ósq������<.���8^>"|��sL�i�˺0�qX�Tø�P �U}hתW�/�vѕ����-C��8�y�͢zr!/��aS{� A9�����M?t�r���`����+�T�Rm�086�'��8Pq���t�O�J�tH�ԫ����٢���7-yPkk�3PeW[�#���0^�ߋ��ȸ�;sRp:�U�5wn�hv�tM��Rj�i4�-�A\h���ȇ��( ~��Ӛv��	�¥�&N�3���@��i��vi���	whŋs�˿<�(^�!A(�Ϫ��5;9q�����窼І��ՠ=���W4�7?��^���"WK�|�������O�����FE�����`'7�<�$nɔx�h��,0�Qw�]q>G0�i"]����N�t#�<"��q�l\�q0�W~�d|�����z���L ����X>{F�ӱ��w��*V�߈���bHw��M�
2���9�]�%��C�����ݏu[�jr�!v�	�ǬhF����?e�n���\.r���b�!��H<�A���i<~�ۭ?��Omd�g�CZ�|m�;:�eX�۱�1�p�.�H�o���+��w�._�1���Vy�Ǿ.n���׾��o>bL��}Z�X��B��R&B���HC�(O�<G��|Ԟ�KVuSxo��F�����/�/���I���|{j_��GbzFF��������E<���^]�Iq�*~vePvD�#����o�k�Wq��wb���U�d���QY�6�h�x��*�7![���k} ��ԕ��8m�U�· ���_�CpE���ɗ>��N���W�x��*��?�0�o��E�/����'qR�ܙ��5��tibL��~@�5�|��r��"�>�x`B@�z%'P_^�N`P��Af��ؑ+��o��Gy�>�'ƾo�~A�'k�K�#���2� �Y�<$�\�9����2؊/�O�py�zK؄9�e�d|^: tK/�'����{P_-���q$u��P����^��'�6� �۷oZ!z˨��X�aF|�e�~[C���� ��ʜ@)+��AZ�$�?�փ� |� �p�/��������?� BD��d�tu5>R`r�=��2h$"��+4�A6�πWʓ.�e�k| �^� �ɯ��T�9曔��!|oy04��*���x��~���]�W׬s�$w){?��_��<�ո����z�����ںF��X�v9^x���p����ν���W������,/�-a @�ѽ;q��/�����㳑�d�0y��dP����y��\u�j"������z���v9y�hu��ǃz�o��4ls�}�*�����n�q�����x���cii�{=�<�G]l''yԗ�
aVV�A��\�<ӹ�(߆�R����҉��$͉���<&�e�����Ԡɜ�1nlr��N�(#W�W,�>2�`\|�+42�1��,E\���0����b|��6��}(�uQɀ}d($�y\���������{��>&��br��#J��ECk���8���տ��8��ѕ�w���ì�ц��Ї
��?�Uէ��M%[��6�������C]�?4���.�C<^2�P���j�$��i����T?� 	�{%���N���/��^{5&O��a�7o��O��i�qx�'^$��1�T4s���?��3:�ԗ������]@<�J�M���벐4�8 �]&����&o�8��Xpѯ��*z���-�i�%��2K�+��>[�*�h%=A]���W�R���?�?�P�a����F#l�Ɵ�A\ʫ2�g�Aa4,�>t��]a^�U\_ɳ��T�V�9]���A ���O��5ݪI�����+@\�+:�1��X�D<:
�Rz&H�yяˠ�G�45����MQ%'�P��	�8�J��+L֒V~�E�j|�s6\x�.]�W /䳜� �< ?�}1@�ZQ{X���~#��M~�@���L#�]��+�JG�K]:��d�1z$<��9��ʏ�p�����${̑����W��`�T��Ɨ��Q<���֤?�2��P/&9>��!��p{'�4َ���\0�*�#@t}���X��g3�yS��&�����+��]=�< �yDG�n�)�Q���+]Pi����6!��:'���N�o��~�Y�!�����ნ}����AYu�WғfD��[���ҨU�|O@���N]��`������{�~/�t	��Z�aF�0)�?�Z�nt�x_��y��F�[����Ɓ_�A=����QtY����}��8y�t[���0.>��۷���'��7�ފ�[7�xm%&TOj���6��9w&N��N\�뿌�kW�H��Q�9kH���hG�x���P-e�H0��ilt-'8�m�<��A5�꟯�A6O��"3�����d���cU�z��r��C8��d-��hK��t�14=���sl����ᐰ��y�V�U���oJ7�5�����plt�ȣ~��d{�H��>E��
�����F:�U<1��S} ��o��do�Φ�2��'2i�5�B��[�g\�zQ6��+��^#c�H���u�W]pyC����鈮��h��e����+W0X��~ +aaև�}�����#�|j,�� J�$���<�O)�;�PQ�Jo�����8y���$B<@��irE�l⊮-�����Y6���%yH�ٱՑZe���$��먤��q����Jc�J�gp��䋟rHg�o�Ju�-�N����j���vb"��V�X�#������9�@�JF5�@��S��[���G��A�*�+~ȏ;sd�^q^��_��x��b�Ĳ7�<Y�/���b������~g�z�I��ʐ���+��cb��)�~�F����;��[��f.]�S/��c�4���8�s�:��GV�'�m#W���)9��|��dH��r�_��59�x��u���^��Ƞ�>�J5�������(߾x�g4�����Ȑ����`<�z1�(�[�����D�ɣ��EVè?����W~����1��$��#+��'�c6�F�rc�Lm���+6�^|�%�c��e*�<T~�C^����^,/����ŘUއw��-���_x��x�~3/Ɓ&�=�7/7� C?��������sC�{5�e�',AY��U#��#:�1�G����|ކ�vd刬I��X:4���gu!C�=�':G;a8^U$��'��9�����+�{��0M�J���i��*$��M�7��g?�ǔNv�g�L���G?��(���B�d
���XX��)�_�y���"��4^p�.�ⅼ�q:~t1�������t���<��m�`>�G�{��c��G��p̫\�;](�� ��U>��	̣�^Сr�M��� ����w�a�d'���獢T*�&���ك���l���~w�	�J�awr�!��ήE�A�r�Q�*���-�Iy)|���d:�dVr&���<���qI<i���k��h��:;�((��=Z)V�0��e�� �x��������@X�lD���� àK����C�Lr�If�^^�΢�G��-$Iz�Qg��|S0�-�|�3!��C�oE�"����Dc���~��|���]w�A��<9T�[��y�t8OV��翋G_~����#9��a���k��N���fbU��^�l�zk���~|�n�� �T��8�ƫ�&�o������p$�"V��߾�y�iݣ�֩4��{Jo��QM_a��3O�r��%�HY#��1�ś��s�~,j��x��-c��i�ύ�@�,*�[AI$��Nu�Ρ�$��<��=Y]�!���n𨔗8�&7is��XLO�x���9GJ�爄�mNaǰ�� C��-V��͍�XrLjȌ�82��߻2�vw�q���x������kq����Р}���N�m4��C���ho+����V�O�ũ�_�����'�\R�҆�iO������m�qMO�n�'Q��p�R���7���ɨ���ӏ��7��CVР���Q_#HZ4c`��RwDW��a��� b\�e��A齂�@�_E�Ę��.����J�#��\O�$��E��[qĻ~��Vc4�RO���T7�!V�� �^`,�ǬtB�>A ��@�Ix��%��F��;�Gr2re|�(p=ďe��8�s�Wp��3�ఒ�qM8���M��'��2�.�)�P.�,�B�X�G��Ј&�b�����mVp >�O]�=��J�c`^Tf��)�?wx�0�/7�ځ!��G><r��+�JkJ[w���?+��'��`����v�V�$�4��?᷸o��3IM�F�l=ʯ2����`ZD)���g��30f�0��XT���3�)ʰN��@^�COU�
��B�ʯ6D{St[!^���s��?�9�0Y1(�f"$?�&
u�x9�(��zy�N>�k��o�
N�	B�a@gB>�@�����'��1���L<��s#�Ǜj���4�MN���r�/.xP>��·�y���芑���=����q����ڏ?�so�#|Oh���K�kL��k�{��n{��\Δ�#�kn�U�(���pn~����+W���0�<
(~�n�+<�䒭�4p�k�S��o�>w��=3�j+�,;-��!����<;j'���+ �m��-��b�����^��GL�y\yp���}�ŗ�I�7�����Z�b���{��ԄW\x����K�ƻ�ŕ�߈��c#[F����W�b9�7�rd�q)7bMC�=]��K�^�g�n�*/۲��}��1[|��qG��m�+��9{���V�O_S���GA���!�ܞޕ�\�JZ�c���u8���&�$W���I}��1-���hI|�id�1Fy�#e�L>t �i�̛4�(%c��K�R�S|pE.���5y@Y@Up��FA/�~Y��Ⲥ�Z)�>T9��,GF"�=�Γ�Q���(�K^�
�d�}��9�`%LqS������Ǐ=��t�<h`)���6��v�#�ҡy=�Տr
z8��+\���4
z�\Z�i���E�w��{4uU�/�
`2�C���_����xć�|�ڜ��W�%?��Ɛ�����D�Օ;<&��)>S�a��U4tj���du�<9�doP����H�`��K��k#���F,S@��P��<�G�҃���`?��z����w��ob}�Qv̎i`Cc�ѕ�wu�0�0_�W^�'O��<:����4�2�\��h>G�����|\��uFF��U�I�K����s-���ii��u��Y���ɜ��v� �~���0���)�L�2���h��x�zR�������^z��#�����w���xe%�&���-7>Bea��1��_�ĉ�̱In����ܾ�3�l|�R&C����-O��٘�U��x^��;��ğK�����6��y�ݸ����өS'}:8{�ػ�Z}羦�����"�g�2�L,-��[�g/_�a�9!��aC���B�䟺�m�o?���x�O�Pa�A�E[��j�㙮p����:>u�����j�'�cr6���`t$m��^A͛ �\�iAC�!�#ޡ�re�U���Cn_��f�4�*/��/�X���Oʊ|���/qY�RTy��i�%{�Kx\s|+Yo	������uE��c�;7�o$�G� 9&dy��3mOc��`>p���=�[nP�n�1�ʯ+7A��C�uS�[%k4��P�����? #�P��QH>�{�޽\vFٛR[�Ј�К�xd'��QW�_)�E�/�����)�i�W�l���+��P���[�]8�Nï�W\��������xeP^ߥȩ%MuN�������38�����o6�G>߱"+�-ߕ� ����o�_,����"�yo�B9��yG��G>.˺�gڙ/��v�sb���C}$���L^l��u�pi�!�Qi6y���ʣ�#��P�ȡ��! ˗.ŅW_���\���^�ى�x|�a|�������o�N���fb�ʵ���q�wb��Z�����.�3I	�G9�P�����J]��wr<��t�=E\<j�aý�x�1�1ȓ��~�a������� �vN������@�ʫ���-�f�z�qç�677}+�@'&�bOF�͛��ɓ'�ucs+~���ǿ��/srRiAh��gV�a�蜙�s�\Nzg�6W_�������e4]�|����u�P�=f��%����!������z���C��U���	�=���٤!��uD����l��ׇLKG�ڣ�O�r�.|I\����8tF��pu�nqx�����t��:�1��,�9���x��]��<�A��4��%]�Fe�8�p�y�^/'\�Y� ~%��b���A�@7WQIO<�k����rn�h��u�U9�f��e�Ұ���,��N��o�%��o���e�J#�Y����C���K���9<��_n���H/y�)�?wxA@x����P@:�ﺤ^�K����Z��z o�)���8�SJ�ZR�� ��;^(2�[����l����;@蔕4�gGV��9��.׃Pʁ	+�+�	J��\�����Lr M����-��>� �<j`𣣙3�b�1����&�u�.���:}\��y-H�{�L)� �0�u��m�-r�A��=mcSc�9>���q03K׮ƅ7_�+o�g/���͵������������mV[X��]������wߍ�o�S��Ǒ�nKv	���9�w��0J��XO���A���D~�!���t��I�ˆ����7b~�P�X��Ыc��������..\���<U��ڍ֣m9�bO7^�^�CG��6��:S^�s�nܿ_���A���c!�=��_�ژ?���F�J�N��!/xQ�����	� ��U��j�ӧϴo�͈��ƚx���X�H7Q�y?8���lJWǋ��I�m�oXZ����Us�J��g}�/�e'>W�r%��ո	�J�ᚶ��l���
���O�'�d|��Ɍ�MS��O���(�_�S���������z�'O��5�)x�m2-��@�_Q���;���HBU~>�R�yЕO�ѩµ���R���?���g�p3.�J��ꇸ���O�}��ISc7���j>�:�~���@��l�S��-N���M����R�$}��JO��{���'L����d#K1x����x4��j<)�$R�8ڝ���@<��AP �<ҭ|I�a�^A�k�-��z���o#����_���1a������+�gR��A�a�)9�
:���G�9 �!Ġ�Ʊ_��ϸ
3�`�1Pp� IYw��x�ʥC{þ1��j���)\�s9>����bH����u�w�G���I������"وgkht8O��S������u����>����G���77��g_���G���i�F�đ&�}�v�p�t,��r\z�}`��9]:,C�o�1@��:T�L����}Eǃ��3�TJ6\k�0~�� M�Sϩ;��8�taa>N�8a������oz$��9��|�de��p}��1�P�}7���v�?��I_^_�0]��UoOx�	�I�q�JW��pl+^�C�s� ���镵|�������p-@x
\�v-^}�U��b�fh�X��oo�B�r���7���*����#������}�+N����C�A~)w��%%�"~F΅?�/��d�J� }
4���W�Wӓ��i��8��keV�!�>�7�~�~�����ҳ��YT��CǑ_�7m���kѤL���8kA:?7Z�r�H�G��G�v�6e� _�5�'�MFc%��4x4��o�g~�I?o"r3Qm�r�exe�e��S&����O�> ���T��O�+ub�	�I˺c̰�6��A���%�?��<�c%����y�FO�P<Kj���=e�+�?W~�(����5p�@��|�������)O?�q�oq���`���4��;��ʲ����]\�,�_nv2QR�1�L&�ʀI�,��4�$LZɁ�>�t=`�F��7#`dLv�a�k\�g|]m��m�z�uÏ|j��qG�Q@���^�kl�I'��01�ӏc@FmpR>X�N�e	P��ɹ�X8y*�hR>{����ٗq�˯����+1�U>&q�s$��d�'Y�ϝ�3o���z+�_~9���b�;n�:V���+���ށ7�Þ.I�oG"Qȡtغ-�`|9����ҥ|4�D�w�d�����)�T��_2�Ηǅ���o��M��B�'��ih������� &CVN�7�mta|���U:V��G�orb�{RX�c�V_����ΎW�8��5�G����	h'z�=(n���{� {[���S���{�|� ,ꃌ`�h����8W�5�V�[[87�>�`"?nSV�ϔ��M���ڣ��@|A�<ȋ>N�����a�,RC�?E/q���ԧ�QUhM
�˕m�Y(Y6F4��@�җG�ps��A�	d�Y.u�߰e,+ׅ[PA�,'������'���hP|�u���摱}$L�4��)��c�!-�p�E�����)y�|�_���x��������K&E���5^;���e�N�J(?�ʟ����^6�=�`i�r�g��۠�T�}��9�so��T���7�I׻w�ZO���ih�v����T��	����H�2��gN)�:��<e�=��j�o�&t�6 �N��m��3PQN:�S� ��[��?�S)�; �x�R�(�<�с
�)����v~��,!,K*�	�Ɂ6�s���X�;~Ҩ6��C��=\+����	0Q	=ú߾kg�jy������K��H��9g�yd$�@(��j2�3�����;��{�vw��*@r<�9wc���+f�Lz�&#!��W���������^��AhP���8x\[�S��o������Y��Gݘ����i�W����?�կ���GOb��j�3�j���i�>P�xn.o��^#���^,^�'r��t�ϸ���2���������{����!x'HY�'�y�Y�&�v,��8��$s�����)�U8>�CA�:'P.��孴�?��?�,;d8d� �y��4
ǹ��ߋͭM����� GG-ߖ���eF>�43�f�y��K���%�<y�:�����C;_�X�6����Y���/޺O}�r����y��x�����3�	�q��zʖ�M5�W���)m�c��w��~�pz�AyŽ���6���KZA�(��u��	���
�4�5�I��ԥC��S��YG����^x����T'|�v��#�-^�y�cM�5>�;d%�vd�'��&�>�	����:(}���b�<)bI��>���l/�3��+<����ĥ?d��W�� u��\�ԗ,�C�襪���l�҉5&��a�L�R@9�ü�7}��#�:�}�6zk���������c����u'�-�E}2����nd���[�*��o<���4���ѡ�xAu���ƛ���)W|��@��/ �V����������=ו��q�*�8���n�q>Ț��'I����2�Ҏ�~9 ��pVs�Qy�7y���6�zx��� ��/�X�e�t��#~ڢh)�����4�p2�_� ɐ�^Z�S��D���/:���L�'#15"y�۱q�A|��Ob[���&�cM�#r���x�ġH��l���r������;�����/�d�����=T��� 3�Vei��#p��y�Eá�]�o�iW���{����w	�S�IM>�>N �������z���|�����Ɲ;w�چZ��� �3V��g�$'�ݝm��uzz�O%�!/փm�y�����]�����w�nlln��2�Bg¦n4���	�P�֋���h��.  ��IDAT�qi��+���7~
rqa��8FV�ԭD�����KO�+�pT.Lt�i
�a�C+Т�Ѕy4@��
�n�v�A�<�mB8~ϓ��|4�H�&u%4鮻���6�.l'u��+�S���N?�\e���i �i��	�vխ\�%5h�W[z'߼fY ���6������0Ǯr���+i���f��Ŵ��H|l���C��9�Ҡ�9��%͋�Q�Que>��!�?K^k���FA�chʖ�5�`Q}U?@>�y��� ��ɯh����� ����(���@g��;<�#���A���<~[�[^c��$��K2���BƠ���J�*�?p�*��*݁tUnm��ԏ?�2;M"��Lu�_�Nͱ__E����y�����(���C@.�&����ԍ��i��n�
��j`���Dj5�(:LKȾF@}9ѫnu�NW&J��J�GE��^\N�s'U��OLv}V��o16�:�{ü�3 6N�m"��U��0(C�|3�)��N*.��DO�Zko'�7��pw;�����<;53�.ƕw߉�~�����;1�����8fRG��qU�gY\���E���g_�Mӄyš��n13���/�O�/�I��7!�$����{�p|Ӿ����M�=Ɋu8�]��r%̥����=W܇Ů�0/��nа��.Y�$|�L;^�3�`�u;>�x�7ŷڭ����"��0�h�77��s�}�D՗'�C�~��
�/���+-��7߈_��x/���"����r�;|�Q$pTH�NN83m*T�"/;خ��Ϋ��!�*8&��-��T��G=@�W�T��B���� +��V�3@��6�?�k�#u����Z\W�4��ça@��κS6�q^:��7��L��,�tʁɾ�-�>��_�J�����g��h �y���PNy�Җ�V����)���My0�WV@Y��������F��r�R���s�1vx���됾���o��qk��b~��NB.Pw�g��� ?~'�vP[����4OD�����h2���i<OД�(Ihh=kl�����0DҒF�7X�Uw�N�񠛝�����C��4�7'[����jK��;`
����⥜;��<c5��6��H.��k��Nj���&g>����34}��7/§3��|S%���]_�C�L�,T��}tI��y�i%P�S�7��Np�x�}W�\>�Lh���1+�hrDN�V�nm�ۉ1�L����sq�����ę�^���\�+ON�ߑ�I�a��cfhr� T�WNI�	Z�y0�Q���*�!ð����(4y�l�'�l�u���M�̀�c����:��t�`̮�E\���q^OOV��^��$�����̴�ٕ����A�J��v��_͗��E���çj�+#��K[��ǎ�d�C�����6��� @��o~����-;E/�=R۔s��E��n�e�����u�ڔ|ۥ"ذoy�/��]��ǵ'��L$��M�i��e� G�'zo�T�48Ϻ�0����� q�~�Q>�՗�d�\I8Y$1z�<� �G �k�=d>�O�K�o�y�J>�VY�2N�zI#^!�$݂*? �R|ଥ|���[�q�Β߬�Y}�����1/�uY����g��r@٭���}����&m��Ȟ��W��[q��|8~3U8Nd��C����X@���@���?f�Q;a�zڀ8b%޽{7��'���*f°Q�x�tb��V�;������ }��e��1W_�AkW�2x��,༡� zH�|u04~�`�ק�:TZ���25�
�t�I��2N�.<�S��|.�����oډSgB�uL�#>skZ�i*˼�	Y��/5 UqB��r����+�w��>.A�W��H7��i�T�q�IƉD+9���=[��̦ǒ�TU�!�鉘��Q}r�4 ��cdj&f�_�o���~��]X�C�� H;�Fm�ۼl��i笛J�vi&5~�;�Xk=�P�$��[��Pm	����o��p.��h��j��������@�rк]��쒛٩7'I�
�ȗ��'�|���O�,��Yw�%��?�q�p�x�D[q �jwg�7�s�ړ�U;Z�G]���q/��}�A�z�.x���[Ɵ��g��_�Ҏ�^�w��tf�D��'i�6e��2mv q?�	�!N��S�Oۄ�hH7�m�4�<hy�JbY_��� #y��W���A_�5.b�y43��9���y?���ef��:�l\u���G K��6kG��eH^߬V2�2�+��9f8�I�4���C�C_~������-^uCϲ9-�YSV4)�}$^������̎��V�W�ju�G����A�Il��#_:�n��93EJ�87�U�8�e�.�4�86��j'�K:u�,c��E+�?Y�����]$/��X�G����A�h�����/�J�Ը?�7��i�*Cq�ː�d�NsO�Q2��HD���wP!Jz�+o�1h:m�mhx)���7V�VUy
4�IU��U��{�98���`�N�)�3��Mޟ
5Hjp2 3Q�
�u=Y�ά��y���s�
 �ع聉Ni�#[h��&��9��d A��ޠ1�) �ʻ�x'7�U=:�� 請_��"�;Qqt��kT�8j:֤��mD��neH&l.&���v:�����c���{��s/��rHz�!)+E)��y3�d�� �5L-S�E�~z��KP6  �e}&�45Q(�i�,*(}��`�3v�&�Hq�}�S���B7�:7������-���$��ann�m���~)������)�N�R)|Ж���WH�xAwzz�:�q�W��Yx{Y�R᧧�\��KSU�V������ۀ|;�y5E�7ۿ��{���ܗy>6q�J�vF�ȇ��$�94����4ڔth�+�wM�Ʈ�)��cs�I�t�GL�Ȗ�	�O4�� $&v�A��LN��]�c&m�z�'>��t����m�hYu���T�85������`�Zqґ5�ۂ'X�N���7 d�<B�C�Cߖ�:�\�Q� �r,O;<�����J�����FD��Rh������I˺ECu�b��#���LY���	ǻ��-������[t	����b��N�9��2���v-[O:��z��f�xj��ZؙW��+�2z�Q��\��lC��<×�/_1�����A�Q)�z6���9�'쏁�z����+�8zp$�`â��q�7lX 1X�Y��Nq,�T��Xt���G��A�$�@����tT���&py8q')�U�Rt��9�ҩuN����/t��w� 0(��]م�V���:��J�$B���'|#$���)�q��L�?k����u��L�'<;��gg�����vid� F��hT�#��Ky:v�q`匲��NO�B�m�@�8-�/�������o�ʅ�pw�`����rADm�$��]�;]��H#^�"@9�	@��h{e,��,�.���	�aG��1蹇��*ʑƑr�'Ǥ��T��j�~��7�~��������_�k<z�(.]����T�w����y��e,/��������:mZ<1��c9K�1A�0�h1N �j�������� �����d<)=�{��	��hh�F�:�-(n�8���7�� Ǥ�S���2N>���;?����h۝�����OZ)�v$Ǖ6*�vZr�q��e�S\>���="g�D�/����@���t���XxU^��@��Q�������e/��������X�gd��t"S�f���ʀ�ţ����9:B#jk��]J�їC�]~�^��O�niNS�t��C镖��O/��Y���o�*�^g���ZB�b�]��� �B�{!��.��T�Y�?ڐ �e�ChG��3�� �
e����§.�/7�ٮf�ςl��u���H	��o%
F�o������C��i0���2�4��՜�d>e��&_�<��ã����e䊕e"�� e8x,�O��	��;�,���j)ӄ&9p H��<u���F�ΡӤY9yn�4 �aC'?��8_����AT?�*@��h�������  ��]�l#tT�N���a1ۇ�������tr0ha����2�o�w����Й�2�qH��&��zL���	� ������b�b�9�{�F'g�|��@���B̘�(tT���e�O�#��NZ�j�Ϟ�;���'�qfHC����	��8*��ݷӄ��@ͻ�����!NeIϛ������D��!98�{;�����C8y�>��A�'q���_ ����a��<�p����f^��	ʃ|s>7طZ�-G���H�K�<8��^� :���Ui�	�ݓ��N@�"N~�=��{0��N_� �M��ޜ��1@
c	� �c�5T�������jb�O�u�|�Ӆ�����j 9c^����6O��3��w�QJW�/�N}�+�Nî�2 �*�O�R���vҥ��֯"����,�[��;p��W��Gy�ũ��p���R;�N��R"�4���j/�̝�����ߴqt��2�S�>}��r�1H��.գvs)3\_�C�ym��eqC�ji�� � �{C�Ҡs��s�z���s��x��(��S��76ß/���\H}�D�y���	�����W_�f�T��n�d�n��w�(8��Ő���`�@�3�!S�����D��r�	4��c^�F^�0��1�\�怕ԡ�۴s�G<;�=u`u~�2�L: Lb��p=L��zy�gA��e�	k�lB9�0�Ω_q�'��V2�R����`�a��No΁aݔ�E4�c7ƃ���>Rg�䁲�����nU���.�$ߩ�� �!Z�y�;m�~��zH�M�^dR�/Y1!���x~�*�a5�6h�-�E8���-�m����8z�Bə|��L+�ʔ~�*SaX7 ���a��3?|#�����O�Uڰ����mQ�)��&�]/�Ω�U9O��]��m��E �w��	����yNIu�ǂO��-��Cg�������p�p�xj�Ix(ف����9a8}X� G��(��]}�4eM+��$*Ў�@<�p�a�'��vLǦ����3�)�)�۪����M?���JfQ�eҩ	9ޣ<�k�~A)�-L���ĘJwә���!��~#��v�Di^t^6P��K�b�͜����#yi���S�E_阁�}+V��.Ż�ϰ��c������v��it�q?'�s���`(�&u��H�C��*�����i<Չ��,:��1��lqp��N�,�`릅܊#_9a�BH���8y iZh�'�r�}��/ڙ�֥~����G�<xöK �z�R�@C$]�͛7�Ǌe��0�O��g�~��\:a����~��Es9�{��4Yu6�`��_��D���(%z:8݈>m��Ξ�=[/��.�����r���j���&>`�\D���iaz��n#P:�������$�(�sm�IF~�W�t�����F>|%X"�e��@
�-չ)�,(��:q�A�z�_֑u*��&(~�g2#N�aGΗ6$+)ŷ��_�.�L���Fg�8�=���YSs���QY�;�j2�G���/�������dЀ�|�`��:�x�^�ܰ�@�(=/(�J���5!m!y`P%�#������e��7#�޹��y�����)�W��|._�����n�_����W�ܰ�N7�pivow�;^G�C�#���VmM�W._�ٹy�D�99`L�|�yIC�x�y�M N@���s�cC����:���?}N�죊(���v̫��N&�NE�{�fS�ت�dU��#�Sf������	�]�qޤx���i��d�N�GcoǶ�O'��� �䌩�ڌ�8�	Í���	?�W�����L��T� p���_�2�J��m��S���?X��5"'K҈7eND���9B�j{A�#�����4���)"��Q�p_j�0V�~���oB��x=��|ƞćO��_ڄi6Ne��|x8J�A�����|�j<|����tUu�S�{��ċ��[���A��vuN?%G������k��h���,@0ݦN���p�a�<�;a�?��>����1��L2��p0<��2���	��C��v�Lw;)�w���yO��~�� ����L}\�']�L�iM|L�r���Hǜ`���gY\&�%��Sq�]15��dʁ!���#�?�3E��Ф��(�8��s�����Y�]��}::2XT��4� ҇��g�ֹ�Џ�8�8@�5n.O�'ޠ�S��N����7~�h���?�i�P>��u\��t�RR��hO6�vY���tw]Z���2��	��4�SŁ�C��D������A:Ӂ� �*�n)N�Sw9�8d+�+Zq��뼗����r�v�<Յ}���Reځ���]�S�ҋ&7�P��Cϋ,���Mi��ئ,/neBEUVz�J�1Y��H}�ű� ��eȃw��I�!P4)�<v.I3@�|�6�S,L��7�
�pS<�9Q���6��Yq䁡l�Q�v��i�HcGW+�c�t���8Xی%�z�w��8�.��wm�g._��7n���JtD�%:'�ڈ�U���%��h[ґ�~�	�e<C�\>����&) i@����7�QPy E���:v�:3q4�S���F��(��O�y�q�.-�N���29/�����V��3e�-��ϲ��[�2��Ў)+�2��XY�_z��@��7���C�=�<�{��e/ȑ���`��c�����3iֶ�" ,����Iα,���������x饗�5\�0��zJ �Ӿ���ݍ�4
����w��{o�x48���j-MiP.�,�n�lc�g��4�J5����t�F����Gө�.~�m\����H�,O�S��d.JHz�����W��yl�2tjҲ�1��ا�?�KM}>����:᷉��1z�3�l3�Y�3�_���cM6�Y��KZ�N�f�V�H#���G� ��gD�� �G�f; ɸM}�:�� N&g s33�'1���P��E���D��.io�φ������e1B���6<	���~�����t9�J��  �������Rf��N':@�*b|�X�p9��e+�Y`ئ�s��p�pf�K=O��$v�Hl�[�0.�8�qr��)�g�:oXg�cȫz�+���H$�t��8�uW<�E3�ѓb�Y�>d$��"h;4Q�)�@�?�^�Í�&���C���w���c�����~�}���{_���j��[q��J����)T-��U�?��������<6G��yJpp���+��>��Qz�r�iJ����;<(�MM���q�ݿ��*�%���e9����zʺ�C�5VB���U�!�nwp�F��ᶤ}���Rƴ{�Y~.���6D>~��+����ˉw���x}h�P�+>��(�����E������s�=W�|6|�>@=9c����KJ�B_>�@�0�_8?fx���j0��Ż���x�ˀ��4���i`%�N���N�3:'�[�A�i�Љ�3�g2Ȥ��:G�Q���_Y�����+?��$=��Չ��t� �t�� D�@ȱ��d��(��X�n"�Z�5t�DN��"ʹ��k5�y��sJU��������M���.�_�i�_@��s���k�a�c� ��  �R���G���� )�H���ʞp��de��ꇚs�����Uy�gb�-{�z(B���?�/��ѺU�A��(<³ >.ǜ2�l��Ӵ��9��fc���"��LȄ ��y�FF��mд�m]�L$���Q�v���͍�[u9p�Y.$���J��q)�<vѠ]�t��N�@/�ȱ����B���z�z�>�A`��8j�*�2��x�r;�L=�K�TM�?�3҈�6�#�ہ�`����'�4fv��N��rQ��Q+}�Yl}�U,�1�;<�)M�3�V�K��&����8�ucnv.�gg-�����v�(N�Ѽ��΋/ڧ.B�[d��L7i;E�$g3N��g+�$�|�T8�b�Q�ɱ�����X��ۘ�����Ǝ���Ь�� �8�?@��T=�.Yt�����Ű�����+�mf��{��x�`A��9���ܥ���K{��)�բ���}��)����5WL�5c�'�0O�C�gV��	�6O��) ���������s��
�F�qu^���UG�@[ �l�3S����`��!�]`p�C:#����:3�qu.���<;X�7�ȶ]W���1���SPu3��42 �P9Sy�3?:�N��(Tuу>򙠩U�I�&E�r�����Djp��.�����~e+�F��_�B�����O�s�wh��<�N<��PjC����l���*��R)Y���v�ӏR���-�L&�e�J���m�\�·N\/�9
J����+��0������Ư��t��c����d�Ϸt�|ӻ��R�K�y	%/b��Ϗ���Z���~�T���;DV q���岊y�Q_ �N�~�
�����'J��H>���N�g����a0�pSfȌ�)���)wt����=M��ܴQ��'�2���9���&}i����S^���LL�]��[��ݝ���6�	6p��.��N
��t��YY9^�x7�x���)��=���]�z�n��N8Oy�6$����J�\�g�ĳ2�F^^*�s.�8űhE���X���y�9��ztv�����3K�t��������6N���RuW�r^����.��Gx˅�0�g!eJ���i�H�r�p��_6L>q�3ۄp�;D���<�<�,8\�:��CS&xd���u��/S����9w�l�7�?��1PW�����	~�N�l�pj#����#$�$���`�Wa�Mj��Nkh:�ц��Q����
�́�t����]�M=�C=k���i8=�o:/�����?xap܉�zҐƘ�J�F�q��W�yO�q<;T��H�m����� {@N'�%8����	��1O�z��{"*(~+ ���F�J�i�7F�g�S�>U���q3٠T�/��g�zBQnZ���hM�ұ�o��=c`��K���ٰ���w��X���.H��9.�U ������p��^BcJS�ǟ��sE�r��1=�;����@.[P�I�� է�wuDߔ����ǹ�(]Q&!y�4��+}�y"K}�p=��^���i���W��K�R:�r�7�u�2u��SxI�ʓ�d��/��`�扯��4i���K�B/}��W�p~=^}�Q_��<=��N,-�řŅ89j���N���S�q�v��<�����ۏ����`��M�h�c	����-�C�0�[ꂶ%��(�7<�� ~�I���C!h��d}�vV�P����9�}9�����1�x=�WL�*�s�L�������ӌ�*O��������i�O	~���r���~�L�?	�Qf�^*ߤM7��Z�$���e��Ά����.}�#�ǹ�rA>yC��ˤ�ד���\�\Z\�S�@�i��t��y&>����\�7
qNi8�'�X�������T�9#P�)�HT)���F�	$OIӎS�D�fZp�$p��s�����6 h+O���(�x"6<�K��ǯ����2�������yɆ>t.��p����P���JN���5�z7��cS���x�&P��۳����i�CI8��JGMC�S�<�7�8�2OO����pC2M�W\H,�,yrND���~ "�8K~,g�`���A���$� �Y.C���߇W��0N�p}5�>[�S������n�K6�0��C:y�BZ���)I�|M`�G�s��C���\��f  =�����x�n��,?l3@ٽi�ĩ��U7Py���k�?E�h0��A=e�����mҥ=��sr��r��&�+�
��O��G�H�I�	��|���OشC��h����
�f�����=T�bK��n�(��|��ɩ�i��D��儍���(��x%d���%Qx@�=���e�o�<��wbHK��v�
:HrY_�_�N�/�����<�G��C�}�M�o��T�g��-�{��1&Gt|v��S6��354��q{��$p�gv�S��S�t�@g ��o�2�e3�v��A]���38���o��r�q8��7��}�	d�������%<��
ĳx��"�:Ξ=���MYp�[�?�iI7m��}�?f��;a�� �Ơy���~�N�y]>�c��/���aԙ�Y�)�'e�$����(�/��S�`P�4�ݙl9��"��~��s'm��I9�yǠ���e9'�9���9g@4n�6Fޔ!���U�
L�R��w=�@]t^:5���/��w�����D�dΑm��Lǡ�	�L˺�ȷ��)��C骛�%؆۾�<�2�5�S��+��hX�:159T��Q�5iC�џ�M�m�e��>$��$1UPa������D�T�$/��D^�i����rT�.�u��s`�:�-�+�H�F�� ����%��}]|�1ۓE�iL�(���Pr�>�I�?��V�ҹ]��9;�H*y��a��<P'F��)�0 %@L��gT|L�|�w5�w�(:���T�����ٖ[f\;Ѳod�G��i���pHޑ��W�U��ԯp�,�g�z�((!�0B�
y��s����\Z�}�1�"�4�+Y&���y������~�n���l��w��;�����`���Ն+/�o��o���[193ۻ��>:�^FbYN�ؤ�nJN��R��Ryx�2����3�/�ҬP>֊,J��ܟ&}JʴP0TA�ݑ��i/ �g尃,Ck���M������g{�V��ޣ�i?��+잜M���t�{�V,]�SK�nks):����EȔu��'O�+v^i�����]Z+��e�ĩG�aYR�&�t�"��iHΫN�q�,*.��[���g2�M�S���զ��u�;gn����t�Gy���.pS��U�?���ܗ������0�������,I:U�YN�AF�F'Cl����_�smu�%х*�h(���*���'5�9w�d�G�������h�����c��A���]�t���|�~�%p���W?�Q��I�R0�0=�P��!T��^������J��s5��!Z�o��{0��hy�kv�R΁#	�A�}�P�&�Z����}t&^�O�IO=3��D����?�M�iM>��q8�b�g#���@ur7�Y4q�� �ta\��3�s�8߶Ԩiy����5���rB`�7l������"c&P'��:�@E���&�|7�T��uU��^\I�wɕ�֏ڀ6q���JV{)yN�΍�V���M9`r
d���I���W�3ȃ5S�yAa\��_ģ�?��G�cg���o�b�t,��bnV+|��oe+����.�?��dy�cŝ3|�r�dя?�>H~�M���rܳ%	��D>2Nߖ�y܉��Ob�˯���GwO�����)�\��;iK��,�w�r��n\S�+�^������b�e;����ݎ��Q������kWb�����y*��NT��c��mλ�T���#Ȁ}�1���>��Ȇ�pD��P�~�T���
�,��v���˛闧�����4o���u9c#r��ʛo�{���?)Ngf�@�1��)������x��l��6☼d{�V}'eʛ�A/�6N�I��֋~5��0���C��o�%�c+�q��!�49W��5���u�%���>��F>J��6a�`׍�v�S���yK���1�s��X48��a�~JCm����6��Tp��=�8=�<�;�	>P&��$?W:d`8'c�Rz"�� `��t��&�:�;�N�c�N2�g�q�5�Yfh�ȿ�5���?!��<CN^.㲙����I�������C�F�S<r�:^���Ь���It@����t�����9t+8��O�W��i�0pֽȕ�-mg)��E�x��o����|�
����l��܋���I�s%/�g"���HGmGs�d�35\d�vzr�V)��G�O[q�ȡ!@��ۦ�����E�L����53��'�<)� 4=����o�T��M@�*��c�ć�c#8��.����G���mo�Ʒ���C��۹�]�>�{��Ǧ�����m����Y;�"">�6}���AU����-�Wp9���F�/�(��<M#����p<ƥ���ݍ�O���_���n�뜛Ч��bjn&mD�'�v�'rVzm��8�f��:�gWb�� F67c��>�G�}]9q����$_Q��:;7�jD���cTeҿ�?��iW�&;��Ӡ���iOَ�J�Æ�)���AI�-m�n��֥�ȱ��I�`?Z��wwc�� �c�외�޻q靷bG4z#jc�Dc�z�?��e�����I״�����j'�o$n���h���E"[���w��6vL��I�T��C�@/ԛ��Yخ����ҡ���2���A^�-_Ā^��B+g7��R�����+�?��q�o<o���sp�{��/Mg0.��W��H��1��Sw'W�I�˃G�(=kH`���Ńk����2��_�h�!^��Ӑ��
�r9)��Z]ϴ�#��e%s�K��k�)#�֤	>�.�arGVʒfz�ݩ���X:�βN�i�+n^T7G��#�S�!]4q�*�tSt2^��t�Q����t
p��1i���<�+ɴ����=��Àf�U^_?Ci���^G&�I&9�aDQ���L�J5.�'��{��Q�aג|x���i��4ẔIy;:w\��W|�dX����v�~r�o�v"�|P��Yɧ���	��L�5a����8ev�$y�̚<�Ro�URG��i'N��X���?�S�߽��r{3&�c�����ݽ8�ߏ�N˯c�����vsG��t�����?۵�[:�)G�0����9����l��DM���^r2��Ӗ�G��N�g_�Η��	�)���Q��'��˞��ԼdX�~�����ss�1?1�����_~�Ft��S7�rNG�x��z-�\���/IL0��ٖ�I�𨸟@GB��+�K���#Y9��lOqt	0�ȝyl[։r(�0>1�:Gcyv!���{'r,ggfcF��ƻ�g"���Y������x������t���I��\nGwWUu���+�8v�=`3,�y0Y���W��H���3�l�;a�{v����t@��L��Я��O�JJ��m����ۥg�|�yAC�:�/_�x���e���aXh<���|�s�:�H���z�R��	�T9�:��YN����Qg��?�`t���<y7���'i�)!ޔ�o�����N�N#��|����~��d}��>]�gǫ	�:3�ooç�Of���8�P�����j����e:fL��i��D��r���/�3��r :[	C`~�ѓw�Uq��~�ѿ��\W�!O ��#��W8��C�p�1 hcp-��4��P����x�s���h�©vd0�4�ż/C�3�S��m|V�\6ߓ#j��񘝜�d2���r��A_���r5�6Гym���+^	��t(W��,���h�OJu��l��f|��SO 4jRɾ��h�Ę%���J��I��?MX<4@9�yҋ�	���^lݹ���X_#{1*'�X�K�@������.�=�K�,�FOL�/^KV��(CɧH�2��O��������)�s�L���.Y|Z�]�yO�������8��ۘ�;�c9�X�AW�&Զ�|bj2ά��ѣ�q��Ń�(������}��vD��w�ǚ�l޿�
Z��K|�1�������L,��)�4�g$��|�R<�F+�f���Mx����� I���$���RtC�g�Pc��1�A/�nLv�iu}ɚ�ݓ��؈ӭ]���q*�m9��)������s����d�ʥH��83���'&�i�ڥ�?x# �rǞK�)}��A^.>h��)o��*�z��,�`/�~�ғ��KPYV���ǩ�ӫ8�2x��ol�x�1ez:Ξ9��YO�P���ǟ��c��z'���Do	ff�P���� �����e"�ڤ����'M\b@�i`p�c�jH�m��e��7`d�jp���w��.�p����Ά��BNt��Z��ȡ�|ꄎ�nHعP�����O�R&WR��8L�Y&Wt���	�s$K��W?�|𐭯�>廙��< O�Q7�p��<�O�Au>��_u�S񂪛
Qo�%=�(OZ^>K���
�붏[4�<P�> �J*=�80@�������54��𩜮?~?����a;�N��b����[}�Zt�I��|�9��.��Oߠ�A�e��`��Q����8|L����r��~��N>z���a�Ȕ<���}���q�Nt�\v�,+t�$�`� ҏ� ���+��qAȤ���ۍ��]߬�ys/��]��a�'fbtf:�"�E�Kޒ�`�'2%�08��Re�r�(���@�L��?ʗ.F{r�76c�o����ە�)�l��m�O���o\��s�|��ڧ_���_��g_�eM���q������׷�����;�~Tџ���鹸v�J����w��m|�ŧ"ff��}VA	8b��梨/5�;L�NL�=�O�d��>�@����8���z�|��N��uJ�Voo'����W_E��Ь��;l���1u��0x�6�"y��O��4pƀ�n�M������@�v��H~�ѥ_��7�#�ʱ&�3�ȭtʔfp��{�Q�Ř����f9g����ƣ���gۓ룟��׼O���T�0`�8�f�Iʿ����s��X��	#Ѐ8`�@m|j�ܥ�<����W���̪�O�̎��iR�;�!¹�Wp�΍��2�a�,�7����9�,�@)�h&.y��@�w�4@p�*>�:"y%wU�APQv
��yyJ*����̕:N�|ܓ��=0*ݓ�XaU��e-9h6t�Mm��}�NG?�|�z�S}�;o��������$2$S�;��FYA2Jy O���u���`{v%<����у���������	\��sB���&;9jV�^�H��:̎ə�d���������7�w��x�����G��woǔ&��gWby~΃+��k�<=�Dܚ���)��S��%�g�]�޳���_銧=��#m��9�Ä�RN�0aYO��'Y&�V�_pҍQ����Z����O:BW+��ׯi�=�SS�V��B[Η�1�7:*�9nw��=�����Ԏ��с/� �@ʄ,�n�+�F�����j۔Wz�TW��24��V�ȁ��~��;�~GF{s3�'Fc�׊�K��;��ŗ_��s+�Gld{7:G������bVtz����?�hɁG�n[z�IxrjZ���6vdO�c�޽�Y[����Egm3*��I�f�8��-&�뼝��F|�l�7?@��G�����Wr���i�l�񉗒�0���y�0v�Wc��!��'�n����������1�0���C��AȢs6��V����lnx����*���|~�R��y�<N}���C,X��*�6T5KVӗ��c��= ����g��
�+;���n���r�U�����T^6������!�z\���S�?Fx�wª�p4xJ�fR��jO���7Yy��h���&�~t����YH'R�|�lw�]u������`'Z���������������q:`�� � ��<��,'My�'<��)�jR��)���txe @���Lg�N�p�+�j�|
shH��W�`P+]X6�,��\YOS^ib��M��, ^��=H���'#��"�+�H��G�Cu���!r����.���͢���Q�5HV��];'\>V�w��7�����a|��6n��h=z����/����D{{#�֞h�\�^���^��Xl�[�Q��Wժ�ڦ��Q�VЕF�K��=�S~�K{��jw ���K 0Y;�*��0�>IG>�O�;������L��q,��sMœ1��?]�Dsla>fΝ��/�/��N��|9����sp�B��t\lO�L���|����)X��k��?%��ٗR���Y����[�^:��K��Q%$����Y�RfxW�aI��N��bO����8�޶�L-��K���� ��_��X���qa|{?�8b[[1�S��?cj�c9_�r`FԆ��ӗ�%É�����8Q9.[����N��ƹ+W|�y��F:�o\$�d��Ű�Hޝ�u���Q��p2�V>P��P�|*o�x�D���s+Kq�U��qZ��Q�������8+��� ��d�8W�Pf'��G[z�k��{�욀�qw̟maĻ_܎�h#g�r�����e��:7�F-�I��ds���	f�,�Yf��x�b��N�!���c�(�Z��s.^��<�dB�Y���,PW�_�y��z'��0�{Z��Qhgs�s��W������Щ�\Ɲ�I��L��{�H*��1m���x���(K�;^����Oj�d����\�����y2-s�Τ�H�͗Z�%�L]��4�[;a@�S�y�E�8[L���kޕ���wHAw��ʫK�Цv.ԄggG �<Io:EO���1����*� ��~�k톎R�Oj)����<r�w'��uJ �-W�V��W�:�t�N\.�p��Ȁ���|�w:�r�����ލ����ی�n+f�Ή�:��֑��;<R���w�N�'z�/��xM �P� � �m��`��_G}�Ԣ�*i�L e�I;��ew��Ӥ�s0?93*w�d5�|�M|���q"Gdyv.�,,��1�8�;�ȫ;|>9������q�&�N/��֣���{z2&�b�꥘9�{�T�m�>�Fb�qۚL���Y��MZB��<�8ayN�I7�R������ؤwB��a���w�ź��M�8	�p ���c�����n��Do]N�����#Q5�0v���-�'fbR�׸ƉI�5����seK��.�{�N5���#�7��#q�_��޻F�+@D�X>�t�y);�k��
�:gqr,G�+{��r����XXX��>jGk_��-�1���qE�@G�s� {DǮ�jt�ɱ�tx��7���r����s�c��(�$�iy��&�rZ�U�
 �B< {d~��k�P�JF����=��~�'��Os����\�e��3e<YP/%㳲�N@��y��	�#F����'W��42*o��ذw���}�1ѡ��e<6d2�U7�Ӊ螂�S�����w��� :�O���7���Ɏ�ĥ�ʫ3�y@�q�H��JH?x$�M'5�Ä����I�� ;+�lԙ�(]����.yP)zt�v��x�� tB��~ݩ���c�� G��v,sR;� �<���c 2O�A��6�r#�#���P]� ��v�W�W����K�(�I������ (@׿�S��ݶ�\��t��f�4eT|�AYAs�w�Z���,Y�Y�������S�\rc����9'���	�άhZ�gx�*���]�y�D�����۔K��L��N�hRG�K:T��;�JpB>�	8��f^y���x�����w���Q�d����_���ޘ<U������;����钍���L����޶��ѢeQN��K1w�l��|�����wh��ο���Ё�����.J�r��s����5x�� �TE	қs,���T�0>��W�����V쭮ٙı���t���K�qI�k����c��rJ�9g�d��:95���ӣN�N��^d;���G��iKt*����i���T̮��S9n�����)ܗ-M�\iK9~�����OHg�&�2�>��_h<���1�����?s6�eG�+����+o��_x�N6���Ң���ð0��<r���v����\�t:h�����8��ĮH� N� dt[u�i#�C�>�˾�C9��P$����jJ�+"ȗ�9`gcQ���q�/���d���<�s�Ѹ�D���\�ъ�'����6�t��]�@F����� �U������#����S��= �2�~9�!G&���'	��a��@F\�A
�䓍9�����P�Z>ݗ��@P��u�U:�&�xQe�5�rêˈ6��ĳ��av6����%p�|5q��\��cp"�n8yy�L���A�t�����ӯ/)��Z�U���yIp9L��]�5�._�#[�(��A���8!��c(|B�^�h���Wz�S�#���ն�c��#n���9�=�n@�؊�_^#q���O�t[m�7�J�gϟ��rj��9���7�2+�.Y8˕��w�j��ā=�yPo�k�i�	�';�v�dE	b��{�p���Ͼ���՘S��on���'165�	w9ϭHN�U�9&�w�ţ?|{OV�֭�t��ވ�{������\��i��ӛ���g���k�|���zaׂ�`׀~X6�ԑdh�1�ocb�6J�mJ�r�cWH9�����~@g�p?Q|�T��G�pI�+g����ݽ8�;�#�q�-^���`�]����������N����v�hM�~nj&n�p#.]�m.=�5a�D>�C��}^$Ɇ�]��ߋ��d��Ř�#v"~��EC�ﾧBȖ�e:6ҷ�K�"��>�S��|^�����0�i�5=��yL���h���I���œÃ8���q�ڵ�T��&�v��;�,rhS?��.Ҷݞ�Z y����5qH��\_�S�ӥ�}}4e9���qlg�4n�6����km�}��Se�Y��|�6|���4�\�b{G&ʹq�L(]�3�<�s�VF	И<�\�a���!r��)��P�v���e)�ZE/q�q<
�I<h��ay�/<��:��40��D�<���^�n��LP��L���UySG�$O%ěA���ٝI���z�@��ܝY�2�t5�C�N;�I�J����2d���jxN~�3�Q�n��c��	�ɦ�N̳do�x�	YO���v2�����0�ԕI�aC���3F���g�g}�Nʖe2n܆Px�G����n�뜀Z�76�� �x�77��z����Ӫ��<?�Ilvv6�T�	�Y��e��H�ʴ'Q�|�d�q*<)�l�� v�`w��,c�5����k�F��r�8/���N��/���iT���h�P=|�Ew��3wcJ���Z�Sp�i����і^x:t�o�ч���?|;����^��w��_��0�q��:Ƥ�iM�_x1�\�[��S��C�����\ngx���ѷ��E> ���������@>5.�����8"gcLN�%j����s�1K�ً�=��?�����O>��/��ӭ�|-΅(p�wZ6uV����\n�D�%��w"�w#ox�SXje���8�b,�ܣ�s1�r�ܸݦ��1�a�%���}��F�`�W�^���7�K�P��]�-\>�����DN�<�yW=�POm7�)ˋ1+}��X�x.��W��	�25����19cv�����u���N�x�]�
����׋�����
���1��Py/��Sm]s��* �}��$�鰥?��Щyb�v�r$�1�T6��T4@��Ox���9<����qc8tO����Ӥ:�t�4`���M�N��35:�#=� �Xu�$Ԕ��C�Uc�.�V�0�!�(�l�d�&����0�� ���[|�B�n|���S��)�Ny�F4�dY�ծŃg#���w.K�Jv`�U6�.0��0if��Ut�Iz���
`׿��YՖ�g�˴f�qvC�]J�O����Q��1އ��۟[�`���cF�X�(�UrnvZ�V��'�����{K�:fpb�Q���3�4� 8�]냉Be��"�/��/x�NR~��2p�p2�~,���>*>&�xG�7��tcZ�.�|��o��������4�ub~��M�-���&͛�pvq%��_���7�܋7c��r���p/Nڭ�b�U_����y�/Ǹ&R��ny� ��^�3�Ϲ�=��� A9n?r4Q`��L�ś��+P��*�#��ҞdTu���h9�}�;w��	{�뫲�V�K��陸���q�ͷbli)��H�>xO>�*���&F��c�ۑ��w��ؼ�]��vc�H:�h'c1'�Wy̳��݊-��󯿋���X^Y�����"^p'�A̲��`#ȡ�m���=� �&��l��G�������ڀ/$H��G�NK�S9er$Z�����?-G���JW�s/ש/M��>��fD�K�{��A�<�E�N�&[�;�K���C����n���_��o�����Ǥ�ȷ=��?:�Q��l��_�cWK�K�����7j����dW��;� l�.�F?�ATF"�!U��13��t�R���b�p_��/W�z�,3��U��;���?�o!������9���7�T�,�� ����E	�F} '<p�%9�Wǜ?4n�V)�\h\�R�,�Y,�n��b_����Kiv�x�Xz�U#
��Չ+��h��H
M�?�|Po�2%>����0����=a���u�იҀ�L�`�$�2�`Ӟt�l��� r��	�pl���9� ���d#�OB�ð����:rRj��Dg���2��$Z�3妓�Y�'��ǳ��+:��#�����a���k@p9(8�����i�7WMT�f
���nz��*\��h�)��)d�؜Ꜽ�OS�Lp�>�~Ji舎&�Í��>~hl��?��g_�������ai��� �KIg�bbi��=M��鸄b`V�����;��s�Ӯ�72"6@�u�,Ҙ �p�Ҕ7l��J�6�,�E��W��=88��
J�� [��X���}ےyr�4�f�͊���n��7��_��̟]����М��at�w�`m5䮹��$7�	�&�E��$�QX:\�oK���tޓC��rH�$�Li��#@^9i ;��W9��A8�V��(��-�_}���[r��?��\�c9r�V.^�k��g^z14Ѳ�;�q��������v�Ȗ:������J޶�v鎝�IM>v�e7��ٸw'����5�u/&�sn�ǹ����F�a*�7��qN��N�D�#��t�m���i(�g�/�5�I��2���م�Xo��k�˔��]�ςE����$�
����b��O!�r���ӑ]t?=!��ك<0^z������_�"���N,޸�ͱڊ.#�Uz"[�)C��.*�I��(�ƽ��6'�����|��3&^<f�^.t�D��^���"T���>�~v�bni�7�����%�c�1�c�0���+����i���S�5����.�~�#3�C�oH����B{`΃��KY��`w���M�1^{���l󝿬!ڼ�vV2N._���C ��� T��������ŏ��{�����dHkkk9�#��)�|��e"��M=J�o�1d�:V}v��sxC�[`�B���L�u���T��̝�2�r�Fq��<w��x�L����}n�
��¯�;L�P�T@}:/57�+�|��:�^���9)�yK2_�>oT����p��Hp��4���Jc"����x��Ѻ� �����ۋ�'�c����|�$��D�Iwtj"�XNF�k�''�S���CL*̞��wF)��9��ƾ��1IS@�C4j�(H��Qs)�۹tpR:`�4:��Ň_8��1M�_}�/oǶ�ѣt&�Ŭ���N<0s���F<���hooǂ�^����rF�<^���C_�?jK���%��3gblyQN�&�@���) ������y7�OC�I�ѳ���a8TY~8������"�W��6��5	w�����v�NO[��1��s�.����[�"Mz�89����ǫ��}�����f� S���,�x�E.*F�������Vt�Z������r����eR��U���,����.<.!+|T[��m
������.f���j-䣻n����ιLw��ٸ�����@x;�l��PxT>��N5�Eϯ&aBg��n8L8��5>��Fqʢeb*���#���q3��x#�_��ssѕ3х�t��O^�uU_��I��. y��vR6���oN���_e>��ό.|�q��[,p��_�i�9Ƣ��d�o�����_q�9��i���\	Ѕx�GUg�e�?h�#� ep�H��������
����Ⱥ	��r�k�}�#� ���/m͋@�&�2��c<��.`�:u�������~��]�*|�U����#<�;a�G�@��{�����$fE�ۀeaaM@�)Q$l���X!�#Ch���V�%�Bu�iP$14��2�Њ|�>P4�����#礻�(JO��K
�=ŏ({���M��Q����9y��� -;�V�I�2(ӡ�.���.���Ї������A�"��~.sd��AW?��#��*��Ԍ������[݈��협6#�eQ��x���8�#�ք��iy�z|b:Z']MXj#lEm��M6ܜ�6���c�)��e��Q,��ɓ~���m!�Y��9�ޱ����a���������x���"b7&x�{�m&1�eQ������Y_��/���>�0v܉�C9�Vt�Wh���hmm�J�����#s�|�\�$m�����,p�w�?��/�:�y֎����ec�S�*�G+���q�VJ�6��~8K����0��VcwsU��d�Q�|노�⍘�����~�Ɂ���������5r.;���5���]#\�֑'P;�NM�p��y�1��fzf6����p�%>`O����;�α�Qr7i}q������7�{�z����q�y�լ�W�~+�W�b�h7��lǆ�_p+�1ۨl@G[92�=h��������6�f1:9-�oɹ��v%���Wq���c��8_����A 0~rY�U�І%r:S�G�s�H�<;aN��\�?xL{�4j�o�7G�'�i�πC���X,/�zz�xe��՘؞��U�tp�	z�+y�|�y�4/����x�eU.	�>�+p�4
��<� �*|q�"�[.t�C:�J����u�K�g�z��4\-=#/�,��0�>u����~�����{�h���21������#'�����iH�4��W��~b�U�'���eS���ʲ!��y��Xe��N'�q<h�NV����[���ȁ4;l��(���$����G�!0�cY�W��:oN ��gC�2��:9z�A��.[q�ֶ=��zRZ�Μ-���"�h�dK�>H�3�	�o$����'q�d-F4)�kR��c�:�i��&Pہp��¹�1:=�]'� =h����1)���J� ��ǡ�YZ�Bv��8�nʂN��È�s�����Bq��%�	M�'r,��܏�;wb���1#:\��N=llv6�oވq��y:p]����?�ͯ��QM������Z��{뢳�d5:{��(�;�ĕ��Lo����V�ߋ���X^Z�ٹY۶��G�I8���)��N��`��x��a�:�I��_F4ȂG�JJ?8���|(onr*F:���ފ]�;��_9��>]9	|�p^��������ؽsW��폧���gvv�;
R�mǘ]���`Zz��L��15��F�Z�^��׬t4�:N��-�����Jy�;��"�?��=x@�<:>RF1%t����P�8��8�0o�n���[7��_�g.]t�q-Rp��$;��j��]m��	Y��j
��1x�K}yR4#v�?z�L����q�~K/܊��N�&tltV���Ы��J�V4�Qj������ �b�'���?��XI����4�"&����u�rʀ���ӈ�#�9�[l_ eM�I�N��C*YG���8\��0�M��I�R@cvA����� ����f��U���:T��m瑡E���6���yK�о�E<Ӫ�?��Ш�(���~;aÍH��X��v-O-�˧���<q�0�S�1髌���xL�@�sW��D��5���8_i�R�����00��X�S�E����e:� ���x:ki� �;hE����I�&;�@+�I<:-�����1٥.:9��o�f9�����7q0K^���d�e�)i���x��&=?-�¨��&�ə阙��%�ݭ�����'K:<-xԒàU�aK#�V�S3~c�¹O¼1�T�\`Ï�c:p�|�Qɫe@���AZ��DSmB&�� a�H��a���:��DK!"�6���q9����8x�0v��D�9arr6�/]�K��3�/��>�����h-��������N�w��p{/��v�+G�3^Jʧm�����3�	zx�~���;s��)OY�n.ڄ�(�1Q��T#g�Pck��8�lP��Pg����%�����{��4���S9ɪ�F�� ��t�*��}o�?�#GsDɎ�ύϿ���������8��r#r��]������֏>�cޭ�v�X<p�X�Ө�Of�m�;Î�_J;M#3S9���	�O��_���n[��_��N?���ܟ�r��>�OE���D\��s�8�����N,�w|v1n��R��p��y��vl�=��I'Np�w"<�GN=.F��ș��]qIW�.��&_���gW���e��������%���y��a���z��q��Ija��1x��Դ�Uَ�<�*������T���*���E�(M�ù�iUV?k���)j��M�iZ���k�\�3VA�Iƫ�10�s9����Jœ���O�/�B��+%I0���F�M���88'�Tő��#�p���x��-/tu��v$E)���~�/�/Ĺsg��7L���x�8�{����<����75a��u����	e(�qh:i8c�1HA�v��[N�;��/;FS'M��y�F9�A|�ה'�e�crY�I�d��Ɵ3�I����cC/�?|���r~����}T�n�JY��$W|�_r\b�Mh��Es D������>}	L���m���R�����3+��Z9�ɉ�@��<QF��i���Y��/����1�|&��53;#�8�W&�*z����(��%CK�g5q���h{��K3�Tg9���s,��2��,��<O)��M�RFO��� �fŇ�����+T�ֽ��Q�#�1��/#>���w�qYhfn1ξ�B�}�X�yM�A;�E^B�h&�n����w"�ۼ[k$:�����<+�s�`yڱ}�;�:�z�~l���S3�w��͘n�g'ct���!2�m	�����L�H��сm�se�u�t�i�rr�v;(���ػ��'�bo{+F��i�(N��1s�~!��{Ǟ1މ�M��cY�������!��@}<�qt�/�+wrqW'�EvU���+�<��מ���3���:�'�	љ�e��t#�A���R���������r�!`܂�u�9����j��w��`���(q\v��hջ����Dk'm��Z�x�2Zڗ�O����Kq��[v��Hl��_S��sg�m9_o�ݯc�ƕ���U�}ĘA�|�~����~���?š���8�^�ָ*P��!7£O�Ȥ8mk�W�3.@9r���T>����]�.���P+�Y,�;F�#-��'��,HPt�++���9���L�6��6�\x���RY�p�#{��0Yo:2��M�����}q�g�����Xn�t;hqF��\z�ڵ�=b������T��c�N�+<�;a�����C(=i��6��*�N"#�Qx���p4�]�QǚʀT�&�>����#K���g6��W~��$I�3�����sP5���r�+�T����a�)>��
�v��G�����Tw�:$$];q��4KF��48�]�<�
G-��,�Y֫�dM�x��'��x��7��_�{�ə���3��Nm�Zܿ�S=;�6]:{&�]��^1.�x#&����ޡV�Oo�>��2�nZ�k�cǋ{�P��$�U"g�A�?����1�0��
x�\��֝��ZO�F�<)J��U;Yx7��	|�j���uM�q��+	Gq"�VVb���;���o��ǵ�ia���^�6k2��c�	[�-ǄI��y�E�oɗt����G1#�؁<�C�����:�g��*p�LZ�!V�mX;���sRv�9�#��&[ MY#���V�ý�c~�>����� ����uv�hu�Q�9�9�;ҙl�N��9�|~kCN���V��9��ڡK?�^D$�����)o\���{�ŭwގ�W�J�j'1�=P86j8/�/��x/���qП��p��Xʻ�~^H?^�Qz
��K8���T����A��6��O��.�d|ꪫ>��ۅ��d\��x��W�#y�<y�[���d�3W_y9^��;q�ś�lI���}k����}�_}�'�q��c�{K��9S��1F�s#��>��,�,Y�H���5�I�`?yR�8-�GM)���9��cGHzY��
�W*�9��]���p��9���|3�4��AG���q(pNy�i�r���G�٩��e=7�k�I�#���"�z������G|�aG8v���X�n0q�u5@�i��S?:��p�'�I9aeX4��-��X͔bP���8��@.5d�T��F�s'�a����ѓ��ؠ�����嚸�� ��!���a@ǫw��6��|~�$��o��9�c(O�]�;aC�4����(�d r�xT�|��G2)h���k����qL�DOg��j�|w76�|[�yWfZ��̼�+d~K�)N�ʱ2�}`cK�1�0KrP�5ط�v4h��A��0j䌹3K1wvE��vj|ʃ16��^�^�m�U�Sz''!O�Q���i��JKY�3R.��������@�u�]�c^*g�xc3B�8�F�4&�fc��٘���5��Imo���do�����M
`�t�WӒ�K��җh�iR�'�;%�nT�&��qi��)�E7�#����Z�#m��?/T8o��!��Yq�l�.!!�W��=l�z�L�``�QrFm������Ʈ�{��%[���+g�4&Dj��s��ԄW�Z�GOV^]«L�����EBўhp���ۚ�.��f���_ř�7��R�D�S1"Y,����r������}]4iUh��r̈́�S�5�j�&�e���(L=켢7l���{S��t��P��ؖ}l�YE�GKu-_</���<|O�?�-���7^~)���q��U��T�z<���x���œ��>v��*���v���Nr�N��J��Ks1sv>ff��{�������x�����{�� yȂ؜��X3$�~��&�st�bP��!i�ݥ��n���0��L�-	8AФ�Q����5_�#N�gY�W�A����X\�x<jh���#�p�.?L"0>8:�hq)���7��=�8e��}�(�#=�?�&�)p]�a^��2�����a����z]Eu
��!F0��	0�6z�l i7IOG:�?�cL8_�I�8�?�8H��E��#�J�" ����B�&v.h����_���琝�S����"��H8`����	�'��gj���y�L���/'��7�YI����I}(R~N(�޵��^���c��/|<���w+�?eR�O�Lk�bJ�:{1�iE�n����w���23�������j������b|i>�.]���%L�19>��H�L�RN��M3)��QA��Rұ*����)�ԑA(�t+�C��m
hٙ�t�N�9M:�;�|��݊Mx��O���k������{�4Ξ[�w"O�v�᧟�C��`u��FiX��ϸ�)���M0㪛��*v���xɃLGrL��6q�O�I�ӳ�[�<�����zj@��y��q������r0H�>!�K���$���b�I<z����\��/�m9�۱�>���&w�]�NGm����%�k\�^l��!����r>��Q�����˶fn^����8���~3<�E�^c���DR�S��ѻ�����8����*�A�Yb�	*G�FG�~h�7®92��vL�tI���1��������ם��PǬ&�.�������_�B�X|���������"[�ύ7�M9g�^�����?�]|���� H����<Y�=w'G��}e��y?��69Tn���,���7e��҉�$����1��.%7c�{��Kv4[�Uv�!� �	����`;��H�2�����ˬ���Η�̧ Zֽ����M��h�F߮��Ӿ(=� �l��¯t�� � ͲЦ�͛�}�fp]-��4��C�^C��M�F�>�k)�_�v��yϫ�+0͡�ˁ������.Gb�et(���^��S(���2w��x�I��i�ð��e�U�L��t��~�������8���4@,���\�:GGOLM��$U�62̿ y���u�������쨅�|��#`<�͎�|��4�s<32����8�B1�iB@������X�V�� |6ftL��㍭譮Gws+�XYOO�����(���*�}�~7�q����8Z]�'m��-Ƒ&���bqI�{��y	���T,]����D�+�K.D���f�X���v&ѡ�Џ����b�ө��`�����L�����÷�q,�� ���������{��:1Iy9'S�c�?7�������mM�k1r�V���	M�=19gϬ���W�k'��y�(:�� ��V#b��u�K$���I�%y�,������0v'H$æ�&Ic,�щ'"�ƹ㍭6�F \TmQN�`d�9�M��+G�����K/�y]�߈�]ِ~�ʍ�s��1]�@��tg��Cx�őK���䜌ND���ٸ���q坷ble���q�щpp��A�2�e���vc��B埡l$�TN�|��GNu��2��\�c8 C#u��0}��θd���Νw_?<P�ʶ���b���&n����ΝϿ�U9`[�ywtA��܌���9؋�_}��ݍ�ދӝ�8�W��BgBu�J���jy���/@��h�;܏��ɘ\Z�7��o~�!eI�����tώ1�����ʥx�K��b�~�������e�����i��KB-�͇ν8-�)�9nI�����<��s�<}�PG��M�X9�~�Q���9��i�O�R��Ay 8�����zY�	);4��^Y9�r���,PO�#����0 ��Xx"��'5H��0��/�j:���I#I#d8W�x���'�����9�u5�ׁ��#�$h2`C�2�S�Wcԭ�$v�D��	��2�<=� `Yk� ��\���	0�1="�g��!(����2�]_�Fw��"���OON����3�	K������<z��͘nh�b�#���gc�Ƀ��������96�|�jվ��Qt59���ؾ� N5�t��m{u7�	sle!N�mkb����� 61�ȓ�T2.�Ԗ}$CʙG�L��)%�#��4����s`���tH"�'�!2�0ٶ�z:a�iZ6�Ƹ�^r����	�9��ӣ��q�^lib<]ߎY9$�8WLf�����2�N+��wՖ]���/z<��P��N�� U��:s&��\��/��̼'WV�d;B�!����ɴQD8enoǀ�����L�$�����y$��Sr�zf&�#�����_��/\������8=j��ށ�|�AN�9�#�F� \�����sî�G�H�c�+�y����li�E�'�����t�;选v-|��Eɉ�sZ�!��NT:������W������|/����}�i��P��-Hg�Ewb��!(-^</������K�=ދO>�$���8|����X���%�͝�x��Q쮭�8�Tki!�>�1�ը'լ:yK>V���G:�D�^G�׻r�g/^���y���`�|n{�eӦ����TC�;�ݧ�g�O�N�֬�T�*��Y`���7sQ
홙Y�/ҙ�lϻu�e���o�[�q^4����,$�91&��?l�2�'*����>����b���'�I?Ǜt� x�u��ga�Q�h�N����;�B,--f���R���O�=��tª���O?�Q[��9�O�� Y�a���ّ`˕Q���'mt�#��;H��<8|�?�:I����#�Ѷ�`tF;/���pj�y��)�98�A)Z
6���᭠�~�_T���3�� c}�>߀���w�۔�D�d�8��q�'�o�����tf�rP��N��	��L	�ps-�މ���8��'�F�Η^5f/_������Z��;���wc���r�6����~;w���C9X����H��ˤ����sq*�����X���8�ێ��c|��\��=���"��]I�\�UC|��7�C��0�[^+����n��̈́�����w��x����bL-/�1�i6В�{Ўi���+y1!���Y���xR�:|���N���1����D/8r�"/��#��H�x.�_���{'�����-yp�W5)LE��-��S�iZ܎�ڠ`B�.ގt�M�<lAL�juN�����#!&n�+/kS>��e�$�Q'f�XP��+�+�q���x���Wފ��/ǓG��Z�0���7;GvN�c�33���F�z����N�v���I�ǣq '��[o��_��/\����=���Tvo�~<��e|��D��ø|��A|���Q������˾�;�ݰ�w�bC:�Ar3�f���2T,�����J���!n�/'�1� ��zr"�u�.�?�06�.]�.��Ÿ��;*;�}��$�n?��A��c'V�-����3'�w���$���#�R[up�:&���@�!��Hlj!���'_��~����ZH!��Y�F��̤���W��B��΍��˪�~���9�
c��x����´Ǭ�}]��M�1h��x�4��\��	B۱�s����/�+�]9xP��Ux�'N����3o�����H�>GxA����q;�:�cz�|25�p�b�R?�r��՘Ԝ	oU��d�!H6������?9'�Ƶ���1\���N�	��a�W�co��Nr狡-i�!��W9�hV�>/�^M�n�oe��å	N��uγu��L�7��B: ��j�s�T&'���ND�m0Ӥ����M�z���H���e'��9"�f&5��F�V>�O�0�aP^�w��[�׎�{wb��w1à*G�oB�6u�L�j"����f����q��sm2�����59jX��� �}-�]?Q���'�UY.av<1Ok�_�N�i��ץ�6�JT�:U�^�l`�j���,WHv��}�('�q�ܻ�̀Nȃ~��	��E�x���܂&����:߼��9^#��Λo��˷0����4�)�'��;9L���=s�k�;=��|=^��/��k�����?Z}��7��f��+�ǎ}SG����+>x鮟��l�a� n�p�\�7'.�p�(,S����P��Ը��;��w��w>�¯��|�(zrV�吴;�GNz���������x��7�W%�dY�=�C�w �vr*�o\�k��_{1�ϟ�iM��;�Ѿ''�����g���7��ַ�cbK�����Ņ8s�t!���/Cu�K��86�6�"L�����R'�� =8I��:(���&.���"0�d��)��ͱ�w����i��+��̋�D�4�u������򻐧m�|Ee��lUq���)�m,'Gޟ�G�L�J��"��=�&ν�F����C\z��ӂ8��b99٦�y��5ޘ�&�2[��3�y9(û��%Ƿ�W*���2��T:b�q�XHqnNG��Fq�p��6m��iZ��	(�:�:Uf��>]�8`�@.�CWU�s�
 i5�p�K��������X�b�T��?	�Ǣ]ǟ�$w�0�jdv��ݻ�2@��#��#c��i�5F�y�ձĩt����^��T���i�(i�|wxh68�4`����0��x�T�C�ס�&���^����*g��S��p^���D�lj��%W��� #u��aH���f�͸V�J?�d9������x��tT���J,^�3����b�ۋ��V<Z��;�bD+t��Q���>�7��$2��*������I�7�i��Xȸ�Iavy%���|_K�dA?�7���I'W��$��@`0�	D#J���gi��C�2�\q΅:�O9ʠ�Hrl��ģ�'�K_M��dB�w�`_�%]�\��i!����?v,�o�'<>l|�֭x��W�z3N��娎���c9�����Cg�����"ٙ\���a� �@w��Gk��bб=��<
���&�S�;�s�rT}om-�����ǟFowϻ�8|�|O6�'���+/Ļ��x�՗�@��7��c�yD��t�b�|�x���c�̒i=|��}~�a�����ݻ�[ی���ky��'w�T��윿��g��`X��k�G�?�C�B�F6�M{��C:[R���9tЇ���J�Ic����i|��Ö��p}=Z�G�G~��؈�'��w�Mˉd�gO}�Pŏ�'�+�����֎��(��E��˾� ��Oƚldg~*�����������7^���3q(�}��f:�t '�I���~^��)�}�
��~�n�[%rGl��8�'N}8'<́��P���xN/�,�o�V�31�B���a�2�@�#�o˜�WZ�C�xZ�>op�x5H�r��XF�<|�юfS�(3���?f��9a���Ccs�� �����{pذe��� M �2}��Ȱ��KM:2pN�ꟃ��<*"��=;E��cM�w��|���Q��*�8��e�j��tO�J4������#������\
��NC�E�sҵ�Sz�@�λ"�Y���A��r�/m���)+>���v=Y��������o��,Ǭ&�3�������q'׶�h}+�V��)t�ز(�o��w.��6���^���O�4q�Fg���X:>�]��K�<1�S�"n��雉��>ܾ�Ѿ������BVD����F��l1
:I�1a4&F�crn>&�c\��	�������)��.ou?��b�O�U?�U=)��/�H?r/���1:5��wr�|�x��Xz�誮�&���l^�
��ĥ�T�\R�l<M	�ԇ��C�v
-M�(�p��T^��d��9���%���^T'�\����>k�<=��G���qt��.FB�X��I��ޛ����W_���񱜪���c��N���T�z��x�������b������%���Gq��w���h?yS�'��iv�T_[����y��l��|tŢ/�[l���G��{r�~�@��q�a������,��!����� J;������E���m�EI����X������h�l��(��!?G�/��q5n��F\�3��
�veo�q������ؔ��m9|+�q�o���%Ϋ���A��%Z݄�����CB����a5�!m�}�1ܴ���ɫKyiky�@����<i5�&lY�Ь:3='q�K�<MN�>��N�\�9��-�N��G��Sh[�8�Gǡ����>���af5���9���=t��
H/��M;,//ǹs���g�ǡ�S��� -@ҿNXG�����6Bu0w.� ##��r�	�A�1����z���Ss�\ˀ�L�r����qB�A~��v�tt���Nƛ)�)�A�S�M�r�')E?�!](���td�����ȯbyo$�&��Kt[r�\A1őSzr�0d9*q]�4��qde>-�aL+����b�ރ����2���|,,����L�h�8���nl�Q;X���ꛞ��3�.�/���2t[q*�k�7��A�ɡ��沑F,��0{
[�L;"23;���5뚁X
�>20��
n�T�i�|�:B�����<}�DE\��)�'�9��XH/m������n���,�r�[9#�4���%+�|9A��\^�-�a�eo���Hu�5�/\���y'f�^�F�qO���5i�Dl�EOa�伞HW��X�xg�Wm��!��T����� i���:�
=�`��Q��*We��R)O�2�if�Y��K�nĴ�|J�w��fkb4.��Z��?�&.˱X[{_~��X��n�Čd�����t>��H������<�����^�l����~��r����)(��	P����8������x/�ڍ RF,G��hޱt)Y�5�&�)�4rr��|�Ў��5��2�ac,>N'R7$��rc>ѳ������v�b����5='r�/��b����g���ߤ���w�܎��m�Q;��#9z�glR�y�Wy�.���Y��_b�W�Duعq��w/ dJ�'��R���9�P3�Κri�m`&6yؑ�Փ~���O:�e[�t���2.+ܺ�B}v�2P�>���v�,P����p�2����3G_ ��U�1 6��#<A(_��Bo�I�r�J�nҡY<�^yU�i`�?E��^���1P��^���fC��8'Z��RU��Y��A�5 $J�e`��NƧ�e�/��σi�_<����$=dѿ�s������@����$3��Q��ᓖ|'�d������2>�[q
ת�.m�X�����r&}.���S�*�2o��e������$�դ6*灏&�l�6���ʜ&���n�mm�2Sku-:O�c����V~w�З��'��}.��Ay���=)�ʙ����'#1�J\�&O�OSQ~gO�o����v8s��?�L��D߻#@O�	T�c�3e-�9�FV�w�&v m7u����ESW��Z%�M0�x���ӍJ���y�ҥ�r�/��4hH���f���>7v�p�x���l�Դס��C���ko�g_z)F�:�m�3
|ʨ-�o~�u<��X���ؗ��f���b��7�r�qu9�5�D�U�Y�w��P�l����#�_������8�|�QD\Ư�n��Qѻ��+����:�z���Z]�/>�(��y�Jg���w��ˆ�yJ����2�}�U<\��u㼑���e��v�t�O���jGU�M�{�vl�џ>w&�V��#�H�V�qC>�L�����+��ì��+`'�������;J/�����O�α�п�'�X�Oq�SŔ����hK���)?	����u�|�M��Ѯ�Z�~�ѿŶ�ҽ�]-�T�e�O1{�3}�z���!^�������@6��bl|�2Iq����"eV���M֕qr�t3��%�̨%��<b��/m�#yຟ5u�=����t��s���	�,�X�pt�څ4]�w�5ωG`���Z�3'po�{�����$;����Ȣ�H�-�\�vH��q��8O|A�l~~�9�.�U���}��?T�y������1.V������N��hd��Z0?��2Z���v������D�+��Ƀb���lؤѹe���g9 sՔ�N_�K�L�����7I+���8��i��S6�ܛN���7�W�ڙG�`F=�G���� ,��r��8�G�~R��2:�]`'E�u�i��9BZ���!�xO�^W���Q<Y���cLD�t�h{+�ay����ڽv8�X�����h�/��Zߌ��=߀�%I.ŵ%v�T+@�9�}O�J�Ɓ��\�+7o��e95|[у�@�@�Q�+�6�8I� ���A�:�d���A$=�׀��������N�4
C�&7�#����w�=�����w�PN���'�4>��9�@Nԑ<�ѹ����t���q^�>�۷�/����_�[r�/J~�P�$��6b��۱������c��O}��@M����r�,.x�GuB΢87�v�$� P� ^z�-6�.�s��?�L�4
����D�B���-:W래����v�0�S۾�˟������/��_�������vLQ�\�i9���!�?�-��l�c�'���ǜ��r>i�Tѱ�&H���ݐf�hz2�_�9���2)��Tml�4�/��޶�4S���t�.9S7px� ��É�ʭ ��a7��&$�(_�gRF�c�Vߚ]^����b|~1����ヿ��xU�@�z�����������8X}Sr�FؕՂ���ׁ�Ͽ�J\��_��_�U��?G܇4�erլN���u�폏���ǒ�lg����s��� ���<��My�Qi���t�W��X�R��	3�8'��Z���c�~�ӏv�ɇ'����>R꠭i{�ˤ��K��! 7��!ޠKm�P��S���|Ω��Z�-�ڠ`��y9��b�������>p�M(�������'�6����ޞ���z=����sV�et:�W+����Bu��̙�?���ǐ�壋)�(�$�x�NE�s��yM�*�����H��:G9���Z�����qZ3�3�4ej�Ɏ��u6pq|�
fZ�Tz���r����/?�(��Uue��m '��9�G��X��0h����{�15�vd�H�ӝ�8�;4m=~�zR�9#<O��ޣ��������Ih��6���g���F�>���9��^5.��z�^8'��(��в�/�J���}}e 'uW��HsV�Fq�/��!^��:�bS���P}lҙ`vw���۱��I��q���	X�,�8���7���r�n��Bl��y�����٩8w�z^޼q����]߈�_}�>�<�>�,v��6�r�&��.rH����^�Ĝ�y9b8_"�en�7�K�;:�斜��@nQ�ҋ��Fȶ��;�Dڋ��vH��8��r/��K7�ǵ�_���E�`'>����/bls/&d����9�Lq�q�J�hB=�rrbx�w"�s�Bٶ~8f=�zj 9a�'��T��r9�������1.�W��g��b�K"AB��\���ԑ���dGK�դ}�q@O�.�)���,@�^$;u�����+L���٥�p�F\��J����1;1k�ލO����������q��*Yy�ڃ�)i�O&�^�˿x?��콸�W?��˗��=�r���rx���5��7G�cc2�dZꋾ�[�Y�A��F��*ȴ�
}����\}��#HZ����hk,jnl��U�<7��xK��)+�h�Y��}�C��y�v��4��m�C<Gm������ �7�r�ZOm�_��r�vۺ�H3x3=��L&��S���V�ϑ��U><�1a\��@$:������A�v`�D��N���9�z�I:yM$��%��s0��Ҍ�y�@�']�r`�NQ�p�� |O��qG`0����Gw�L���;u�憔h4I���'�?%o�_+�r�/�)�I�I�Q�ᕲ��ę��q)_����5�k���rԞ�i��F���i�����F�r����u=4�OƧ^��p9%G\ROE�#v�F��b������ęW_����7K�KN�V?V��Dԕ:��!���Xț���l�:1^�+/ӥ,�N#۵���J�OB���N�yA�BO�ЩϞ��S�rtr*�|�z&��>x?.\�h��Ͽ�M9b|���,�?�o݌��ߔ���Q<���X���h�݇ObdK��&���+��g�F�v�&�bay�G��s4��N�jA,�?�;M�+�79'��
�ltx� ;qI�	��!z��N�����x���賯��p5F��b���K�q�	�/�Q��)۪�cvJص��)�i5ы)�If��z�=y�}=n���q�ͷb�ҥ8��6o�)NG�s�ہgDB7}���I줂�ie�)=V��eK�ֈ.���}�8C��;�"6��g��H��)����ƣϿ������o��կ���m�V�����G�t��b�������q�o~g�y+�e���t��G�'�4_��m0�[���ߌ�ÒRƒb>8���4��y�AU�fZ��1d?.O���^.\������i�?Y�e�~{H���W ة��|�l�~�I+��E�y�5����-!����T)k�<39�y� ��{��ߔ_� y�q(�Y ��K���
�	Ø���7�˭W�:��\��1W�e�I�L
�;�hk�i�S`���r��ƆM�_C7_KA�ٜ�4~�;��MPp0j2*�$��O�kȝ��/�z5�r"����Gy� �f8�+H`�	k��t�+���
�2������ ���:b��D���V�=9�Ȱ����[�;�t
��QMz|�1F�cZm�E,�U��H���F}���s"9:�_D2�u�_[��ȹ3q��7����Ĺ��s�����,|.�@�/�4M�S�¿�TZ�!���3�� �W��{f�4y8kܟ���J}��~�]+���*��T�+��f�baz*ڇ{�-=�:��N�����/�{��e�?{>�~�M|�����F��v����Y�Ϝ������Ï��g��ރ�����������/v��OOec�ɱ?
<��G1��g�p��LǱd�M��7�����:AO�`����rc'����v�2��3�f��h���L�LV:N��Z�þd⾶�;����]=k[v4:��u|B��"@�����]���\���E_���]���7y-�����]5�ɥ�q��������oƸt>2� ''�J�l�Ed��
��c��ɧ�3IW�O�Sg�&q�-< ��3�$M0������Y���Q��>:񦕬t�w~��x�c�ob^9'r���+�;��fb������wq��w���8�_���O倱o8.i}�),�s�ϩ#m<-���y�Q�iJH�Sn�jїPǄ��p^�XVD6!oXw��e���S]z!���4��x�:���`��%��ڌ@����1�`~�8�<�/�䥥'ݲ�������ٔ�g6,x-��S��O��'�rЫ�S���65�M�6l�n���4����?�4�c���p˸�H����iƤ��O(d��kN< {@��)>���+ԯ������Kg�+)��r�S'��!T=uLHi�@�c�]_�S�+Pڎ�L�l9��M�Й���$�G��䞦1>�;KZ�]�|!���KF<���S��{]&�ү_5��EW�L���������$"������8���q��������Y�l��s�譟�z���<)>���~H[2`�^��\�p�L�=/��j!�S�<D��ʝ(��=_�q��31+'b�{�v7cby�;`o����t�r<�}7������'1��j�܉�������y��D��0z�{q��S�-;_�r�x��\�h��{�K����{����\Lr3��\����o�G�#i^�S�a�<{X/BG'�A��~p�G�&w%��܌��-ޘ�N{�j<�ݺ�0��=���-���}���^�G��q����R\񥸥�(�v������yG=:9��N7vp0^���������*_�!�d>������)A��[Q�t�d%/��N2��,/d�}ʩ��Q@�_C��N�0xB��6ċd��p��d�R���wqj"��~��ݎ���i���-��}�۝���ވW���ǥ�ߎ��75|&}ll*&G��a�W���"�b�l�� .dCFl?[����~�9�Q6������?��Dx�������\�@J{�#�MCC��<ʪ���P|����:��*_c:sV_6˚uX�fL �;�8��8��K�,�=�Μ9+++�/I�.��ņ���r�;�?���@j�a��ǳF�)[�e��+Nk��u�8F��� �;P�`��\$�kp!�O�F��NB�;��
v���б�b����t4
VY&-���^v&�?�M�R	�Ȏ�=�t(/ӈ�  =�+�,@��n�y�c"�=C�{�C23?g.���ʯ߼3S��>����b̌�c&���Ϳ|_M�s�S��R����xbd"eU���՟�y�F\��;q��W�D��Y{��g���>ȡo�#�Z�+�0���9K�' ��$�M��#�A'� +`G��2�h98g����Uv�إ��iC;���h
��9{�LL�Y�3r������[/�������kl?x�r���t�?61�:vv�x�0:�G�:���=��ƻrH��2ȱ���:.w�ZR��5���:\�Z\�ɕe�Ì�2�Oh����-�@ik)߳@��R��s�߳6ŎW��G��A�8�y\�B��`�`�FbY�qAÔ�������ٍC�#�y�ث����f������+����^|������=�ë?z8���~�����q��:����b�ʕ�����i9��WZP�w^��eLkFѫ��	1�e/d�`f�A��_�$�>d����D�}J�'l��'E��S�ҕ:�_�}��K϶�>?-S������%�e��/�-�d'�v�儩�we�j�˿�y����Ĺ���g�d	�����/�1��L"�8`v�D��D=���̴3���>���xEP�e�������*��t���u�'q�?����q2���h*��
���䜝Z���.�pN`�[�$8�p��v���$t��Rq�/� �(�r�͐��R��!��i�c+<YvR4̓������\��S��8a�2�2(�����6t�^1�v1L��xUA�S�_0Y���@�2P��t���@8x�)�dZtt�䋕�W4ɨ���L
�S	ML�:*7�S�y�y��U���%,:�x'�N���e�b������e�L� ��QH���d��nvx�i��Qd���ɗ�4�qO�'~x��ݑJ[S��e�[�sg/h ��	Dx�8?���Q�U�{U&5pS��d�S3q���XXZ��~ۇ�і3��k�/ߊ˿� �iU��A�Xz���u�Q�|�X���X��˘�8��0�T�XW��a����X�rT�72Y����� ���/P�a:��@��jM�􎵘 G��>Y�tt��U��Oǎ�;��dz>��^��/�V.�Ɲ������X���u �]9Z8S��kRlK�92L�
�)1�ҟx�U�Mဌ#ӄo�n���v5�_y).��j,_�����GA��e㥛�ȟ�G�`B�-����7���P��C�=�WA��d��M��O�%���}�G\VT��0'�u����_�����q����@ޕ�u���b����uZ�h[���ġl�#�n��W�����ү~�����%U̍�jC�'�K�F�sk�FVښ��iE>��%����7Ҡ�z���7���+*PUv�����z�Dh2v��șV\t�ٜ��������;<���9��VV�����������7nDofV%���e���3�t�n�:G�/}��x����Y�G6狗�|6�#����+P�oz�3/��9��G�Xlt� ꃖ���&�)%�J}�~5w�O�c�c'� ?�h
�
M�"O@<���!�p�Z��Zv]�.�9x�3���_�7�?ڠp��W]lk�ݳ��/̜={�祋��ߕ�1ۭ�����T�/N� c �a���V��L(�8 2b��|�824:=�5v�@^�xL
�A������
�2F�e$;�R�阤�A�r�F<�8�k� �t:@upa*���Yc�Y�3�K��8�'��#PO����K�D]:��<W�IҹO�+�t\P�e�|:c���=������k�����nl�'����];�L,��	����M��٥����qUN���Vl�m����r��]�[?{/���z,�?+Mm�����|}[���ŗ�u�w�N۝����%> ��!��+�/���0J�ĳ�G?�X�u�� �4��4�ϙj@�2����<'���V.v�I���O������O��P?��6ޠ���6�t·ˏ�5�K����8��Sr�x_Ż`�ٶ*>vZ��S]�7o�͟7�/���V,r��WK���d������:���f2�P� �Ob�e�@�������1?��x~�#��+/݊�e���V� GrF��׿�}|����_���s<""�g��'=�ONĊ��W��7qU��Ai�)D����/G�?�n���\��_�1I�l�#����� ��OB�X��'G&�L�ѱ˒�L������u��=/=�X��}9�k8���qE:z���CL_���^?!)L^󥱍s��6�̪��z�+�p�h's�Ȧ*R�iQ �R��$�p��S.���fL7�}�iB��0��2m��v`,S����mTPmQ��\馝�����1�q��9�=���z,o�5�U\?���s�㐩]<3k��a$�9��mݷVP�`~�9*�c�#�!�~��B���0�
0������?�����!����x�E��ԃF�qӱ0^�ԽT68��YS:��:fu~�)�@_��G�V܃%D �K��r����7��j��Ԝ�;� P֟
��$- �4E��<�����)q���NK::��3�����'N�J����Y�C2 ����z�����D"�O�hŌ����x����?�c��w�f��ү�s<%Goi.�ݸ������#���ݸ��W��s��Tf.����x�?��K�-���w[�
�N�?X�ӽ����H�Y�?���/��~��Xz���.-�V�N��ȉ?\��0H�&�Ai���TzMB��ԝ&4e�]�! �p����#��ݍ���ؓ3�䣏��cdw+:|�FD��p����Ǔj��ɸy�R\^\���^l�sM�G��8js#z/&G�?lš���[��;oť�^�����H"w�
�SS��F�"�U�(~kG����[ő�x�"e�C�8�����6�py�s��&��N�=:';���Ge���cq�����������Z���E��C]=����A������ލ[���8���q25-;_�G��(Έڗ�;��� �hsƔ��Ȼ(Z04*ix�I�g�'�
���]�k����+=8b ��%�=�H�Ș���r��T�#����+sr̤��8V���9��$�v_�ào�8��Nr1F�x�8#��l�ҿ"ݴ'���N��q��i�
2����mQ:�ı[��v<�r�*:��%`񝼧��H[�;�;����M����uHY�N���Y^��2,x��X�"�;�#��S�x� ��¹���"��-^��N`�ҟ��c�~���;�^S��U?z�vR�َY��8�	��O��&��`<ז��lo�ں;�p�Q�l<𘂌C��
�d�22��Ы2�%��/�K�j�@`gI����T�e=fF�lȪ��a	�H��>��8J5H.�#�&�=0�IJW&�0�դ'/�_��W�g@g�w0����8��=�Hk�6xЕ~�ǲ�3}�pK�$7�*�N#G���ڏ8��iK�<9��c���q��bF���΃x g��7c<&����K/�+o�����&��>�4>���#�����{��1�ɗ�z�+�M|��#��N>�<�L����P3tģ8KR�j�t�T^ry��ܴy��l۲��3�r��e�ī���/i�9�	9crƎ��L�m��~���>�q������X�~%^x�x�����rl��G{w?�G��i��0��}�ޑt16=ӯ���y���bli)z�~3?N)7&���f�q���Y��x�g��F6�"T: ^�V9��t^0�WGEҦM8�p�Tytx[�q�Ǘ��/�z�#r�yOݔ�b�8P�wgf�����'��Z��k�D��DW4$�0M��G�h��Փ<Я��G}N�_)�̐X���N ���:H�S_A�ݙ4��˹�B4�N�>?t2�{�d��#�=�#ꐭ��6N�z��Y�	�	�I���`6�=Sz�i�����Ù�चfC��V�e=�@B>A���Dg4����ӆ�� >y���/�5Vڛ��e�
��	�G�'G���xY*}!��Q9H<e9p�X�����b�����������J�@PI�OgR�O�+�>�C0�?�Wi�1�;�Yܟ��	k ��8ʰ0n����ZY�' �c2�1�9�{y�p�S@��:�N�\�6xpc�]4����1T\���C�AeO9�^ףt:���gNi
�8���"�4�!$��|�S�YJ蕖��᪃���|M����t��92��`� �K�ZFؤNMJ^��mٯ��(&.�f�w��;�'�aZ�Ե�q��[q����8�kwsg�p}':rH��Β&�K�.��kw���O>�'_~^ǰ�'�--U�1�ǝ������C���}��K1=3Gm�<��$��(�vF�O�~����2�8����qs��b�7����D��(p{AK���D����ۛ��:���i;^+7��ŗ_���}ۗ'��[���_���ފ��Q��96{�j!���Kq�7��{/fϟ�.Η����r(�	^p��,)����dzJ���{8�V�����&��8�q��i�W飢�.C{o?���������8z�$$�&E�lRm�R���LHo>x7���g�;���H��'����j������ݡ�n�A��?��e/�)wV�c�HIH���A^�������M��H]'�T;G���� ��6��l�2|�z��o�+��u����_����'�L���	Р .$|�{7	�'ل�1y��A�r�P�j�yr�̨��B�6e#�[vZy]Ό�P^W�ҷ��_ʒ�3n�w��DqBO�"���h��-��%P/ދ-%�ǃ~�I�PENd��Jpɫ+5��HN.���n06���!]�S*�d���_��ll2��#+��������w,�ƎHc���/��N����4�(z2W�B9�Ҁ����KR�@�8�`�st�	?�`R�SE�ǫJ�k<�IVsrv�NsY������_�Wu�/� Ss4�7�;�d��v�}���#.����ʀB=9��
җ�c���T��0��a�aЃO9�>v���?�:�jN�|�r0.\8�L`�[�.�x3.��z\{뵘]^����x����~��Gr��ij4�bJ�6>���w���cG�\M8�xG�#�ڐgD���%M�~Tcg/�U�ʵ��ɭ}�ِ��m�y�����2�2֯�(�����v�1u�PWA9#n����W.��ٕ�?���i/�^��o�o��xC����������q������tܓs��/�b�ӋC�}��������������B'����΁J��兮:!L����k����/ �P+��8z�r�c��VΖ�5��\���D��0��dW�Z�qi�+�9��?p���#��l�������_�,�_|1B���Ĵl[VUR�1O��Ƒz/lP?�:��>�Cy5v��2
E�\K�	�����5���4ʑ�J&>tz�q(�ȫ|y���c�	����̎��%�^�F�S�Ľ�&������ţmW�jC��6 l|�f��,��K<d�z�:�2d9*��U,XߢA^�K���@���,�XX��n����B�;;�vb<�y<�4!�m���.!x8ݾ?K|^�+���x,��ʳy`y������,�|+�<�ue�u�W�v0���x_o��;������@���}��'Q:�����=��Ȫ3���q�h#V�3�Ά��Ϊ��_3�:��9$�&����M~`�L
��_#�;���6�\!��)�w+So�UG��Q�~"��TpR��0��ώ�L�ΡM@�`�*����������E�o!ry�G�Y��o^�,��H��-��:�ӵ'���w��?����X�z!&5�=�3���/c���q���VK��&��1�hQ�Q�����}�@�(�͗Һ-��PM��r`d�\��L^��>� ���v�,�ŉ&`p(�O�cO���Ե��Ȝz���193���u:����M}Zo�I>:�N���#�˛��гx���B<���֊��sqqa1�ܹ��o�=6>�:fw��#���/���Վ�������_�<���N��2&F��
?x�ҝZ�:$A��ޤܒ� 0y�܃4��TK���u��D�~�@���/�pl�j�Θꑳ!Ǽ����h}y;����7��1�r�ۛ�����_�W�ƕ�ތ��t>�k�L���xI���_�����[ح�,�D��A��IL���余/�;���U����[@:oiG9)b+�S�t�B����9:���/l_8�$ۡ�F�JM~r����J�_���������q��]�����)�>M�XG�J�ȴ�J=��	;m��Q���EPC���0���Dl>?yF]�'�F?�	�g>������<B]O�oF"��Z�>k㜃����vc�$�qj�EK��<�����q=::r��e��#9w�@9.UB�z�x�0?�ox�|d���@�0}��T��x���' �pfgg����6$۝M�2\��V:��S}����v9���Li�:���W��"��d�K�t~*&�`E�;���'�H�3#^���eL��#���.~�ڵ�eZ�Ã���WST� &�r�"��9����*�U�u+�\�
T�.�Quy_4<�)��:j3��h����o���c����[ێ��V����IV�mHm9{||9��猐�P��yw7Z:���?���B��='��q��7��;oF��jBG�HYl3����|�[���K�h�#k�\�R7��Ƀ�D$ωL�j��>�Q�HeK����13;�~0y|O�����X��ۘ8l��7>W3r���x��t�x��o�k�����k�aP��1�C
Op �3ހ"�#%-ү�$b�	FIa���?�Ko�Wz�- ����q�t�U?��ϱ��}L?>��np��'&=��k"�����c�ڥ��wW��q��[16=�&��)����7G&51bK��K��dް#�����k�W�8��N�������?����4��y�@/��LK��B/u��8Y6iqϖ�E��g���Key�+OϞ"+������Z�iIk�fRx0_8����4x��1ƺ�ܹ�������J>�x�kQIqU��P?c}�We˙ũ�N�ja���1�GQ�YGg,\�-��8�΢eY@N�qڽl�sN�Pzan�>�H|�M��3�v|�
U�iY��y��u�u����8a
dt2{��\�I�N�<�����roA�*F�	O�e:�r`�X�������90�N�K(���:�]"i���ݔ��Z��QI��e~�t����'yH�L��0�5��ϧp�2FoN���
�,4�я ��'Ƙ~�oO�4��/gN��ŏϕo�Z�72L���t����L����z<��������>Z�S�k��Ixd��4��UOD�NʑР
U��2P�Ȃ\rv�x��@a~Ϟ��_�|7�}7��,EKf�aG�xL�`;y��9hr��e�7�"@7Ȇ�X���{�,�!�2L��Y�ԓձ?�=�&�';b�h��X����>�,�������n�t�=p~��S�7���)�r9�����_�*n\���#O�)�"T�#ms��~��;��f�+��߲��g�«#t���tR����3�z�,1羠Dr�7�19��W/��i7��N��_}���W1u���z�j�r�	;o�~� �x�$�FjW���&Mv%����g�I׌	�5��k�i�rBj����+�����G�$wޠ!uB�Ң���Z��!G�\.oo�yq���=��g��!9$gzD��.-��)����,�U�#9<ΐ�D <�������-<<<B��W�t�C?.�F�jR�)B|��LJ��b�W� Xq�Q_2 �B.
��Fg�Ka�&e�~t$��Ze�����c[�h� �L���#���v!�0�$}��q=����F=D_���7�ĉ�Y���t�M��*S�!kʖt�v�k�U W�Q6�.v����76���1�cH�o�6a����p�x�z`�����xaS�f:t�!��y?�_��Ǒ��q�:���}���~�W� Ls���͹[�@uj�8aк=�7�Tq���V���˙i���� ��!G�� -�z��(�GC��(c���]��N���/1��|������Stp�Vc]8\cÛ�:_�'tU�
9����XN��Bzv�c��N�h���7���n颇�a|�X�I��٤~�}�|y�V��c�~���\�j�*'I��CCU��i�mja�f�g嘙�����gC��}>Hɠ�e���t�Ksv��7�w?���W�4;k-6/�3w('�ɚъ� !/r�w�P��u��%�E�?�Coi��3N�������*�^�ˑ����+����Y��c[�����gֺsϪ��Uя���T9<~��q�μ�y���Z���Ku�MXq����U�G��h�n! .��G�b<.��:�rP`����S�p::;Y��o���6�k��5�B�m3󼳻c��=����)ճߌ���#a��h�[v�g��46l�����<栍��NHQW1 �?R��Ϋ�3���~��!K���EaR/ q�Ma��}��zR�;ar>)3�Tg�yt��r8|��t�n��([��g_��3N"��n�Cv�
Kr�����Q82�;^7%�L'?z"C��Ə�4a)�N�:�R�m��^��E�q��y��ǂt���� 9���<��7i�<:$?	��oSRl<��'�A��M�o�����k׮Y��[��G��@F��6H>3<�q�
'3a�	hD�h�2�)jQ��ɓp�hh4\�`ilt�-Sæ�`<�@�|�V�����]�����j���o�	�s����Cb�9��*���E4�;rz:"�����<�mԁ(�2Aqޑ�4�ŵ���.�p�f>2� E|v�0�`d�g xR�u�����"�~��ÌT�Q��}��,��N1�B���:���u�?Z�����C���&쀏.�����}�]�����-Z���tg_�[>���W�S�2���߅3v��w��w�c�׮�prR���l�4�k����Er���5�=w��QO��B�n�Yh�a�=�K�"��4����:��W���ķ���v]yZ���'�ڶ����T� !�����������|h�~�fΜ��w�Q���bv_��|�@	��]"�b�[X�/�@Hy3:�x /i����x�K�J�����h+�r4�G��[ĩD�1��fc��gl�>i%9�U�3f!�����F�V�|�7��(Yy�(��z���a�eЌz�A���A�	]%(��?/u��)*l������霸I����A�E�q��2��GU*��5&�V�A��J��A����u��~�;do�;<	��;J]�>��6 �/A8�mB���![�!��I�Q�Q�c�~�6�ˠ{��C���/��ɩ�e��;��m�:v�	���ϴ��v�6�cw`=K��MrW�@�X?�T�
�l�|rY6�	
��>����zy:s�����@����Y�������m>,XV��ӴGo�j��6^�j|4jڟ�|8Pg��Ʃlѹ0��Q��g�E���#�r�8� �#A�g�t�@�OtVf"�6|��*.����X�<�c<rNRbP�5w�t`_��k����K^t��>i�/:=�/��+)��KT�.�
�w�_��@���t��4<rGY
��Fa�xSr�\�i�e��i��֬ÀY�ZU���K��ԫ����gW.\�uQ���{���a�N;�]���:��s�6s�]x���λV9u�Z��3��g]�xĹ����RV\$@ڰ�1 *�qB��׀�a���M]�N/�;]1嬓ӈ���u�ٰ�.��̌��|��n{8b3S�p�e9�����s]���@�W����j�ѕn�P�w���t<���	����U�1g 6@ɿ�C6�u�(���'mgԞh����^��d0��D��p�=Mu,�Wq��ǅޮ�	V�R3�8�l��wY?�9�Y�Y�>���A�#�Wku9��ɛ��kЃw��P���
��c�)����=�,n�����(��<�/ā�C7�^G�B^�?�<�'�5���ᣠM��EJf�9Y�M���-�2z��/�.k�����o�sY��&]P�됺��L�2��A@��GԠ^$���hqc�v�r�n�O��o:�D��E!�����56�/3N�g!'[=0�I�-�?�ХO@��-�o�6��ơ�V6M9��Um���[Ϊ��;�E�VP?le�G,�?}�L8r^t���<����RO��V8y�[ �Ѐ�(mj���O�+ �FQ���62&a��Gߝ"�̴�7N���ߨ�Rv ߮�Y�1�(��E\�Iaev� �yU�I�2%jpA��aW��+#�w�����~�P�݀�Q+,g	}D�~�Ə8�D���YK}���b�1� !_���p�D��h��A�R��Պ�	�6gX�vh�!�9�.g�pc�V?�i7����19i�/]���l��)��:��O����wlu�u���wl�U�i�qg�a���t���x�]��ګV���x�l�-й,��o���d�73B���u�C'�à10��0���@ڥ���+����M�9�#��1��%K�����ˍ��X(�^6w����>���m}��.��V��|Ū3�6�����	��J=h�XU��|���ȄYf�?0�|�� q�y�������CO m����~"��b���VqJ'^A�́��AI	�9h���F��pĄ����I����x�P��=ZP�¤.A� gׅΉKVh���t�]���u�A@?/7p\�)���+�"��y¨M*�gu=�D�G��Yb�u��P�wtc��8}�]�Q �	��{D�l��ԏr�����!���z�t�v8��)�ȭ��r(����1S��?י�K,��("�A{� ��ew{]�;�7x��j���G �PwQo���[<�#>�.�&Hl�Oep��-/G�g}�t�#���t��?Rt���a,3�Lhǁ�'lqq�Ξ=�v���!ey��7�P.���p���;�Q#�qݻwϾ��K����4^��ޘ:M��D�<ѡ���L?��R-���G9>�ģ�2�4t>��"���v^)~8q��Jt�Dg��`��&��p�e�&���A�>&p����T�M�5q1@��F�ǠR�pǞ�F
�3 �D��1|0Fq7���',e��9T9c5��~���Y�ٺ����L�i�Z�f[���?���o[ou��v75h�/Y�~��vض�V��k/�������؅k/[mv�Z��'c���1�K�A�����p�u�r]qZ	ٽ^��B���#8�[	�6��h� �N��P�V5��q��	�͕�^�>�I�h��?����=_3w��kv��e��Wk�\U>ܰ�@8�j+�!,������v��A�aȓ@�x���X��I�g��<�u��`�`\��6��s�\��$�隳;g��I��'��e�BܜY�lpB��!=��,Bv���~G� Oԛ�S\G=��w�"���������D�)�Q��9B�DO�������%K�g9��П'@���i��_��',���O{	� ����&�p�Ԉ����,d]��a_|T�u�7��U��K��a��%j��h[�p+�#l��p���������I�m�n�?�X��6.o���Fz��O�Q��FߧNe��*�T�7�~+�z��Bo:rMX���w,��uٱ�W��v�Yq��~P�~�� '�k��	�-�������1�	�}���9w�0ss���;��P��IQ��5�g���jq�)�8> (��J?w,��'�2W�Q���Y ��p�4\txd��Q����q~"�Rxy�@������L��o��ߞ����
�$0��x	=ǌ�Z�q�nQ��x�,�<� 7�	��Q�(t��Z��"�K�3��̚����2BG�}{z���䗶��7�[۰���շ�-��zۑJ�_���/�e>������T*Ή*\B�c�/�c&L<�л�B7 �:��!�i�G�՛0�Am��Cv�0ģ�atJ>� M��I}R��:1��'�/ɰ7�Йo#��V��W�m�Զ�\U�.U���D�?��X��xพtI�� ޳��:H�D�XGEL���t����|�d�oc�d%D� �;}�C�3^HK� ���o��ȄG9�W�`y���/�9)<��k�<r/��rS7Js9<�c@�_g��3�+�"��P�,ȷ}ǝ+�Cv�x%�k ��e�/��@���)���$���*-�:QW�	�<���D~�l29�y����P��V�χ���<�m�k�lop �C�+�*�i�8T>#U��e�0��͛�[��K871�lvn�?���������IO�~�ȈN�eQ�~��קδ	��c�1���	��Ox�|�uQ-��G�#����+e�����⒝;w6ڹd��O�t��l��Y��N���٨��D�����������x�S{;�k�A��V�낀w�� �:�X��=�������0��Н�q'�o�變��1���Agw'�Vt<��H',���a����A���R�M���<������c�G��	'����C8���n��bP���t� q�����,]e">ygTDKEb��V��R�uK2�u1��c9�w�<`K��ؑX�"�,��m�XOv�]���l飷�<?g]�S��oJ�KPy�.������!�������ש�Cf�T7� �;U���0z��N(/�c�;{��}�ݴP+<fV�p��Yx�o��7N�c�����7]Ɋ�Bn4��|<�a�|߫T��N gQ8�GDH����:u���3��.b�'����!���u�i�9�x��i�G�Qx�hd���8ƴ5�MK���t��ɫL.3W
z�|��%ֻ�������)>��t��C8�9BG i��2�.��!1�w�T�p��,�ia��F�+�s��<N�^�����m�)/��'@M��#*�K�<�����GK��-ߟ5z�r9it%I��qPN�u�=��>�&A�}��LW��(B����W�{�?ʎvX�����9����. hz]	���
��aA��/��	��&&p�v�D�08�k�t���1mq���>h��_�6����Nʹ�p�����'�� ��;���H�tꓼ)@Z���0�X'�,q6"�l^���/���7X�o�
㐹���Q�J�>������`�02�FUit4�P��0o 8n�O)>�Nf��i��ߍ,�������*=��"u���$�$ 3iqN��z�AgO�f����� �p\gk�/�p����������?Gy/6s�����oo��pB���AVoDn��ۃG�l��C�{��[�VlsѭLئ�����-���]��_�ٷ߲���S/�S�0���;/<�dF�z���~�^Bo�o�1f�6�F�^я�g�v#p|������o荙��W�_K�5���G��h7�Y��������#���=�~��`e^cW�R�K�ղ��h�Q�7#�g�P�,2�3i*"�hky=:��@�1u�z(�G:I�0� i���;焤I�A��4f|]xE���%O蝈 +���D4��u'�G|pN��%´5~��g�>>�1�Z8�Y.�q��۹��O�Q��I���'�3�G���P����h[�4��l�A+�/�\�M���D� ����?R���Al_���5�Jf�\�;-+����s�w`S��M����ݾI}_+�ҏc�$��-(J�y���rST�ՉuV��Qd�tw��,i���b�>��8��5��I����#N���N���2{����|S������w^�6i�0?��)���"x�>~��	�>y�3��ۑ�h@�G���|��5b8etopE�����޳���]R�ӊ�����x�Ua��v.�g�ĳ>���$v*B:�j�#!��H�� �e����2�=V�ܹ�U���x�5DP�:�\��X���q�L�cԡ�t���%�4���?��j�4��D�x��,�iO�EY�[g�۱��޶�����~-�Δ�S˶�����`�ׯ���NN���0��1^�gF(?��n�X�3%�����~�E�z�D8w�u�����0p�5z�(�B�&��Fq�s�����R�W�|Q�]�R��ã�Ƃ⨫Xc%���|�S�ȫ03<8+�Ó;H81�{�D��W�p:*���~�m���G;)�*�ρ�tX�Y@��q��8o�F>��s���B���3z<xN
�B�$g�PD���2K��g���	m���߄EL�W�׵�<��d��T1�$pFiN��@��x�舴�I�yL��)��s�C?���(�s�	+���c� �5ʊ����E�R�Y5��h��=�mm�ӯo�ӛ_ڳ[�؎n�z[��ze�fM�YA�A>���&�u�t���ڣ�ţ<-����,"�ב�B���6-��:�:9 Ză��qh�.����X��$?y��좔�ϯIc�<�] �����3������7~�� ��/�	����N ��q�����͛���C����s7E��@���L��.T��-}!:+j0O8+�iȫkhq0��:!��e ϕ��F<�x!J�h�1 �;A:��3rθ�C�Ŧ;
Y�~~g�qB�x� ��Hݱ� ��9�w��sM@G����.����E��g���*r��w�o�К���u�<��%c�����0���X��2�ݵ������Ƕz�O�ޙ;���v������W��DU��|�CwʢU��'/��u'&u$)�Q�7�$u���C6�O@^"��4�3�z���CQnB>�:֟~�ǵ��Om�7�9��ҫv��l���
^d����O�GzY�[�m���T�3�
V� �# f�yw9���h=���eWf�/=��1��� r�+�
^�-�N#L;�e{^���!+iN�y���s�K��ӡ�x�:(��t8��9��>ЊN��+�t��!��k��p��G��*�hY���,N�����g�w��Sn?�/ʌ�,�O�/�c&,�����/u�q𲅓��}m�☉����|ܦ�\t��j�}R���>��{����۽w���>�͘�.'kϾ�U_�ag^�fS�K�W�.�̹Ic=g�3}�7�U�n��[�8�uoȞ��V���/a���l��Ϸ[��8_u�37%�Q�=t� �q������d=D��#$/�(�I饫�9B�qH@�%�Fn�N�w����%�薖���[�U�n긡�>��Lc�A�
�id��O�(=�$��ďw�|�):��"�ᴳ\q�V�}H�1B�S<���otF�ġ��²(x>�Gg�/ �WR�Zr�Bt��w}*���������<�gיh��P{�@�7+�h9a�G�@~���8?8�ГZ��0�`��bM2�n�mXK��S+v���쥿���\{Ɏ�M����hS���F�"�#H����c8��|x�mpvY�!�B�Fa��Ef���+�:퀸�5��q
~FϡG�G�� x7���ǃ�8 G� x'ׯ<�;`�G�^��<���K�ʊ����4OG6ڌ���$`^gI=@��G��>�r���@�@?���NB��U���8:4�����8]?�W]P�����Z�O("�ya���x�A-b�q�iK���\nS�x?Qo^7�1�c�k/S0�S��O� �Џz�����C)��k�^�?���?��}D�I�6�C�Y�cj�%��	�)�>�;_�%竡ʆ��ڃ_~f�?��6��ʦZm�����siw���;v�:O����`SrDx�RDłh�CWԿx�=%/�3v/��ǟ~�u ��z1��=E�ț�K�Qw��@<��6 �V ������xo�:c�s�V�X2 .�?}괭�,{�������G��C겝��'N���0Vt� v�ԙ���cV)8o�:h�tO��;:��M5��"ݳy�ő��B��� �@b�	c�5?�2i�xY��紝�(�?�.����AQ�>����ͻS�@%y0 �#��_z)dڡ��C��<#I��8\���,��x�;4�T�#�׀�U7�$UY.Q����B��T�vu�=7gW�Ϯ~�{ּx�ڊg��j��w�Є���|�xD>�,*�uH>�)b�`ˑlG���I:K ������s�e���BO�q�/��UP��1�^�K  o:$��P�߱+��vA{@t�Wgo:G�N�c�E�b�P���&���^ꌗ=H�ETvq��:�p����o9�NI���č|����s�q!�C$��fF����G m�Ilfiq!���{��{�Gm{��pd�u���y�i��7��|�{�$��M�чS?
������X~A�Ez�}@WA7�iiQi"���
�+޸��;�J�ρߴQ^�����m~j�f%wwc�6n߲I9!S*����U>]�����ښӝT�[��q����(	����g��m^��^h�^��Ȇ����x���tDH���븍z���9���2)������9a�_5����|���mZ�9��x�m��N�	PnB�i���9��'N�t (@C���Ԥ=z�؟�7y4��H�> 	��O#����[4X��ȁS@~�q���<�H������㭓:��-:&��(����0�>pJg!@����/����1As|� ���|ɠ87�,��gP	8DeTҐ�H�	���vdu>��Gr� ��~pw(�$^e�cVJ�+%�<��C�E[�C����v��+���e[����ϝ���E�5������]��R�t�c��g�;W�s� C�0���縜@�rr�E8�ȃx쐆0�z>ʈQ����<�B|{T�J7Y�;�B����$:@R�z��7DE����e��g3�$[��E<לi[�E�i� ���?��'1�`�,�(�|v�>T�R@S�~W\�.��h(��H�:<�R���=�\�W)��2F �uܸ���}}tyI���IWG��H�~[���i��G�|�S�v�u��)��7�mA(�酞EYG��ͣ�q^05��EI�v�r4�9p�F��~�ڷ2P��3/_Q�h�|
�ި����u;r����ش�>[R`�tٖn�u:�u�d��ϟ��RY'���\����z^\>�Tm�K� �# �?y� .dF^f���!y�>UF�^�G� �.���H�>��"��)�q�iP��aű�~��Cy�Ν�I��}�/�ڨ�6/^)���~g8q��@��f��FWo������;it:y2�N#��� �Y�.��d#���Ddq�.�]8:�#��V�k�0$8 E�����)zT�#=y� ^���pa)G3t`xHޠ5�;�Qa�#]@'��#ԁq��N�i���x�I��(7�8��Yp9>G����ɰ��LQ|����8�l���%y�sO�U��ӧ��0om��\V�2���ys���k��#�5p㘅s���A�Aa��7�������!��I���H��/��t��1-����7뺨o��H5�����,~��t��ن�].��gф��Xدh�3;��/��� =�^�m��^$ /Bȁ~��"���G��Fn�8.i�9aWEa������BR�D�D&�8ЅwV�9ʏ�W�@U�����)�Uq�ę���m}J���G��hfA��֠���qG��>M(vE�"����v�<>DO~�᢫��p$@3t�S���C�#����	|:N�0�����N��~�g~��9f�����n�A�-9a��Q�ZGt�����~�&&6{���}�e�*m����	h�>k�`��u�\�	�OQ?Hp�����E�s��D@�X�Ț���{��5�K=�7%ҿt���PF�4��e�)�RL,�}ȕe������P��<�qd�o�9�_'N�48�;$E�g6��K�xlmn���(l���ј"�N��<���ޑb*���Q��e^bt�\��J�uF����6��@`�6=�4`�,iaH�`�1�eМ~«V|�RwĔ�{��� �:�,h�I��(��t��;q�GxЍ��dƙqYG�E�y���Y�8�<�aM��=��L"��2�44����Az�IF�.������iQ£� \�MA�1��Sp�Ig�uNyS.p�:@��O�cP����B;L=C�i+w��;�>e2��o�+�w��y@N��>�R�Gġ?w4=�B��_;���>�>�ݒ.)��|�vc^v��">�ᆥ�a�K�1}�˕��4���&�W���Uq��BN~Co�Qz��m�KR��?l�H�x�� W�A�8 z q<*$�z��
�Y0ڧ��prּ�IG�踈w�Կ��J��I��-�nǪJ�)o���q��4Ũ�C�v �i��/�.����~�6�C�tpm�v�%�Cv��Ҧ��@�m�@E�=�MOS[�<*��7_��_���--ڌn�����n�g�h��?77g�F�g��/^�Ko�n��y[][������[�^���غ�u��U�LN�H�,�����k$|�y�3��I4<y�О�[�/���e/xB���.�� ?�:ߐL�q�m�z�7��$����3q������T|v;=/�p��%�&��̙0�]��7xJ�G} �g�d8qN�w�'�_46�qػ܄�LN�y�冘�;� :+�� tPeT�T���x���t:4�+8,�Ɓ ��LS>��w#(Z*:0�����/�d��3S��1�q�@���<w�*��\��pB(w��:7<z�V4���b�188
�z��@zt#�|Fy�:�F�p���:���&U�(��tH@�.�б��ƤY��$��eZ]f�d�c0L2�C�P?�e�{f�\Bg`7�������B��ᰄ�>�#��y aړ�wz�d:�P :ts,����{٠M>r t$�:��	=����¢���*?d$�h!�;��T���Z��3h��S]{.��DYJs^j�p��})e)�Q����":�¦�=��Z�k�D�B��@3��)W �^/%�>[��J�y��ӑ�C�Q])J:���m�tv�LǱ�<,�4�)?���rD�'j<�]�Zu�o�rS��P��#/�֬��ݾ(��:�`�!����٪�ܺe;_ݴ��������z;���ް��}�mNM	S��+7m:� �Y�m3���ip���)��}��
�4�#L�x��}gߍx?�<��6g@���,-�e�&��v˞}�}�?�7۸��]X���r��k�n�U��������6��E��r��.���̌�T_�[��ޖ�U�8q;��Y9mӧϫ8^��FeOkuձx��명C�uъ�NG��_�nЇ�#:Ʊ">u�9�L=�t�.|�P:�ǡ��7h mD���=帼ᜃ	i8`�C�߇<�r���a�Hx1>�Ⱥ�甃�~?8q���pl@�Q�u��w���7��P��l�8��7���|:��@��'Dc�����Ggˎ�{_ƀ���֓��Rgp���BF�:��ػ3à_�� �I�p��S�?�Ʌ�Eq)��܁�G�;s���D�1�q���p>K  >������F~�
:E�	�Ri���	���M� �5!^a�!?>�K��7ߢM��_0ʟ��x�0���N�a�G܉Sv8�J
9]��`:��3@8��N����.��,�a���r��SΤ�����1)e����-��>ބ��[�6Ǉ�U-�j�>pR�yB�T0�\��Η�7r�4j�F8�9�r�!:�-��~���G��FՅ߀�-E�x� XMe��ݟ��~�������V�m��b�O׬��e������fæf����=�cS�M;���!��T���*��.���;���B�]DBqM0h�lg�!m '!�'8MɄn�L������{`[�����[��+k�o��5-Ǫ6?g�	�#�	9�rf���M���87c�Wm�.:��5UnukӺ��Z[��?�-^��8�*�Y�o@����dVJjW�+��5���� �N*3��k�fMr�0�S	��MI��� @�m-��;�c��u�olПtD^hsÉ�H'.tu����z¦R�U�v�Z�~H��O栌ߕ�	<'N��lj�y�bG>o�!G��Dc�����J�������r�dg�`���D�:��y�1�a�:|�����4����9F hw��)������1( �$�L��([�&>:.�	/���N�w�:3����<�C5���rz�k�K�H'/ �r�m�g�Oh)C�F���\��Ű�[�ᅺ���ׄI#��(mX����/�Z����Ad��gn�e�i)��G������1������"b�t��N=����}���u���'3�49Q��$��`<�f�^�MT�-3��4ԗz�E�zCo���	�Ώ��������,�����|�[`\F+n<�����ma��
u�$^p�Yx���[8x8)� U�v��g�������t�hum���};�۷.�2���P���҂�5H�d?�GΞz�*���|g�Oބ#\ґ%�6���`${�1�F�'?m���pri���#9�;��L�7�����}��@S�^��s+R��9lMݐ�}���������S�-M5��2�?�ΣG����w�?��S]���Ɇ�-����5�މ}�)^c_F�y]�<���>�<,Wp�U7�t�<��)ݔ3��nPr#?���!C�t����~zݮ�� ��ys���w!�m(��2a�\���ua<ք��6������	��p���ƇĀc��
������رu��54Z��KR�4��/�u�5�I��A���"�N8�>j�E���ߨ*x9.C��Z?���Ha���C� ���3�����1���e���5?�>h�A�8��~�V^p$'�R.��EF���s�%@0gz2=!��3��������q�dz1@���E������ �� ���H?�+ʊ��^h�>���?�-^�G�>�]Ϝ}�,�޲g�T������ �"8�"�<q�0��G�K�"O�Y�U9
�蠋x�/��倕�����G��*�,T��D��Џ�KP������K��-f��O�p|�N]O���u���9�:�:ғ�B� ���<LU
s�������Q��\̂��:ŗ�̖*�Rm�ml����V��qiw������|��o���w}����r6��l��oMfb�ҩST��$P��>�����Q��s����#=�y�Q��v�&
[�0�4�(��!�������>�ғ���Ȱ�v1���峧�)��W��ʾ�?l{�Xoc�Zk���ڴ�{���O?���m�g�ToT�e�gW��ԙ3�=h[�u`9��z��+aC�+����:D/d���N������h��x"�4�1���t���{~�&]�q�m�������#��A��A�ԩS��̞`Qy���Q^ y�n������p��!=G4o�����P>��������NX:7����EI=��( ����tn��1du��������o</�K-�� ���`�r|���4)wL�G�3�����c�Fz9h�ٹ�&���#�~#�0D�y�F�p�>�����H�Hd�|����$.� <z�=���?&���#�F��#���=���\�#�^Сߍ��Nk�w�����Td"-x����� �\�
sd�����/�_�S��Lt�wp#����	��j�]z��������D��~T�m�ٝ�-��Z	�C��TE��H�F'?F̷1K�N76b:xV�.�ά����8t��K��S�K0�
�6�]�b��6r1h���^q���*�����Kl,�#CpxKw�I��hr3��p�-�}[�ޔ̡K��`�^����k�D�jM٥r]�t�;��!��3�T��t
��r��CF%����������"£�A[*t��(]:�#�G�}[��k{�ӟ[��]�i��T�Tr��]��}[8s�g���6��?��Z7���Ѫ�vv����=��S[��K��I���u�l���d�i�f��Moj돟؃۷mwk�7枞��kp��i�^���8��J
�E:��p�>R�pУMq��N{Gn��*�C�C~�*��gϳ�s�� oH�8�o_�|�y�rc|)���@�I���9y�8`<|��8ad�����$��	d춶���;����xn�ը�k�q��~u0�Q���Lau�P�GĀ=!px�J�;��H�':v��� �NN	EQ~$ntV"���_�Ig%x�+��F��
0��4@ѹÈ;��}q�pH���'�4`�����9_�t��[:%��q>��8Ï���]xI�q��
��p�X�_�K!��.s����]| ����2��C# -��[��/!�-t��C�g,}� ��p�)����������tE��M����EI�{�Zyq�,g���a�,�>��vn}c�w��ޣ'�����ms���h �W�#(���i��R<2���A9�UeHb��SB�����S
d��m�r��ǥzZ:a8V8���쏻|@��r��/)��V�ȩ�v��ً!o��,|�NU�5��l������z[�*y݉?<�m���,�;o=�?_��QYi�E�s]��&�#+��y�r�9���8������g�i
+�����c�w�سO?��ΞM��l���E��Ջv�ߵ�S��-��ޓg����V�޵j�c�AO�m���M�;rH�,�jS��15i+��mcu��>��'O}��S+65;k�\m��5t�u�[�:�6|���j���"{|a��6;�[ȋ]	���iq�
��F���;z;~"�g�\����hl�x�?��� e�×u�<$?������-�	��p���1�`u��K��7����w�A��T�����ع;:�`r:N��	��˅��P�ǀ&�\\g>7�\��%� �(;�t��3.���".�� ( *hE�= ee�&.���c��I��K�F�#�1��O�8��E8�~�u���2�9�p�t@(��ै�CB�Dݎ�C��i).�y�d�;j⠚��;p@4���,p�7p���)�����?d(�a�<�4��?���4��9r�a�@w��3�t¥r5f4һN�C��~�v����=���=��S{�o��OW���i{J�Ux�ɪ����}�4�6kUbi�r]7�w�TN�Y�WZ>�<�M�#��X.Ǩ��\��%�׭f��贝��U,���#��'>*���*�����W7���oK�ʪ\0/���d-�!�\d��Y[�z�V^~ɮ����g̒���7o,����㙫��Ѱ������3�Y i\^ڗ�U�q!��#�=�^ȝ@ܱ�نw���Y�a9�>�):<d��a�e7����U;=�n���<o�?z�f^{��+��iS|U�l��}<[�������������۳J��󯫽�c������S�����v��:��|ϯ,[e~F|Iq������C�: ?�Q�����xq#>%�.?'��l��Y�h܄�G0F�+�J���]��Չ��S#tP5<����g�<��1�u�@8��BƏ�i��]�����	�#¨Y7\u8^�f���9��߳�����_�Ѕ�*:��;��yM��큢�,�A�;4��HŐ�qj��@gk�E�����/B~@"��s�Q�9Ң�xSv �q�॑�\�</�͚/2:V8�Y>;Bg8hg�B~�=�">�k�L���}y`�QIyƍ8�n��x@<��+� ���>�-bH�u%^o�����Y�Y������;�/8��n��i�) ���n�<��s�Y"_�c\�G�	�8�
��)����F<�G*ڪ_�l||gG���1�`������چ[�VC/,���9�� ��e�^�g%��gm�Λnj7�h����`�۫�fѶ�>��B���8>q�W�[�RO�'�x�t�F9�K�/[ki��	O���>�;��~���_mG���%_���F	�v��2X����]`}ԩ%�ON��ܬ�9���-���.I'=�L�f�ߐ�"'�+>D���W���c�xG��˽�.t�,!���8�}5��HK'��u[�8�;5�w4������][��P�}d�A�7h�/�Z���K�1�	���>|h��wmU7�]�	��1�Q��r�j��0�c��֞��=+��?��^_�T�vUn}q٦؅_ܔ�w�Tf��9cب�����m�>�pY.�  �IDAT7�Ȅ��*�KW�ϺFt���^sn���H=c#E�⻹a�9w��6�!r ϟ��3qa�~;Pf�(z逝�N��+���):�w5b:꜌ oMr��4>K:F ����3):븁sj~.;�g׎/�A�$:�2�Lz����d�3jD�t�r�Mb#=つ�<���A�; �����XG�L<�#�g�̟aU��h4=/�aH�HA� �@x�� -ҡ<dYr���,Q�_���8N�HF��<(x�j�.�t݁"�����K#��|r�l����K٢.�W��!-�8g<�qA/�otBݎ�H�Q<��+^ԶY�ƚ�	ɭV!��A/�@eJ}��@{{�J��>;�{$Q�ݞU���@�mͅ9��c�#�2��9���C��G8ͤ)N4���^=� ��q�4=��y9.��NN��'��H/W_n`c�#���n8L2��{`۷n���3��d���Ң5g&�Q�:%�v������k	oz~��0l�)ݴ��5�__���J�nʷr��͜9e=1S+���GB\� ~3���C��k�M�L�&\,�c
R^ċ���(� �vD��?�X�P��}�fOn�1��r����Ľ�9#'l���z�k��Y�G�m��}��-Ιn<٢�u,�&��1<N��o(ǽ���,�8���R��j��QT�Ⱆ�q"K�Q;cֵ''�g�����#C�A��/��xÚ7(�~0x໎�m4�6�xoO�1�AsOqu9r}9���)��I��3g����x��J��0�)����|8q������%:��¬�`���k뮊icp�H����@�3Aċ��9���q�G���$���J�(MhH�I����s���%��p���5�<������ɋ�Ѡ���L��س&�M�r">���!tN3XY>wv��:��<�{8o��� �O8x���(�r��#Ɇ��?�!!q3_�u�+^��R�rg��	]{8���X�>Rn���e����r�xe�ȗ|QL��I3y��#�Lܬ���2�A���QN�k������G{�8��nS��YHz}�\f&����UC}jav֪����]�m�|��P���G��Y���a�j����W�r\��̼�ǟ�u�(�w@�#�2Pw �E���M�qq�.uv =�s��͂h�����_���[V[߲�{f��Q��tSr�����Ͱ���̚���Xg}S�+�4=c��-{��u6��P8�rʘj��\x�U[�r��*׿J ^���#6��Hi�_
Q��l_@�ڌd��+�E_\�v����IZ�W��ń��Ê`�h�9i�����3��b�\g_N��V{m�?�޳5ۻ{ߝף��U%6�13c��^��7n�M�}{
6t-��Y�ͨ�(	���t��޾�Y�WV�����At�$քW��Ó���iw�b{�l'!��H2��%�\c���a����Z?����%'��A�������)}y���>�!c,��_^�c O�1�>�=�8a���]N�ud��F���ff�}�xoo/�w��h\өh�y�����A�U�;3�O�.��lG�4����8�q#q""�L\����̅���Z��s�ah�3���w+�����ᜳ#B�Ӂ X@���� �|y�����^�?)�'uJ\B�!��S�i@ā��6p��x�������p�����K<\���;�$C����R���e`��F@���Y�_��m�t�odq~=�q~�9��{>�W`Tf��Q�DBa�Wb�	ݤ��hI�>w�8=�c�b[�kղ�LMi��3��ٓg���?j;���Q$[.	�--��6��$O���3��7.������p�Wт_�k�E;�s�xT`�H+ꙃ�}u ��xe/����h��m|s۶t��7���ΰo����m�c�%���;]{$g��Of_~m�]�o�j���'�l��=km���ewPUf�fg^�nG3S�ٞ��k�V��¼���^�8��R�A�Yq��l�r�C���9�U��G�="?��K�z(%A����Fӆ;{������mB�iI�fg���>~h��u��؎6w�&']w�r�dk�U��[����rڷmO�{����}�V�E�$-�b�6����';�f3˶r��M-.�@x��M��Ʀ�� ���p���oyFF���C��*�� �O����Fl��Eģ�� {�S7�a7�|�w~�V|}y�����u��د�;��N��?"���A�8�Z�zVw���Gk��|�����Xѹ 'S8p�p)*���*���Ub���e����T�1c�D����@R� F^��E#�0n�0$e�T����D"�����9sM~h�
y2�x^�H�|A?�	��t3*�+�����4��"o��	� �P28\�5Ѕt���U?"c�����	���X�Ż�v��i��u��mZE�vC�Yz"|�X�o�A�?�DY�,����l�����%�e��B���z:vB����x�
�^�hr�
@�>ʇ��sݽ�n��o�������lzzҚ��D��#�I f*�1����>3w���?�ً�����M�[��D�J�n��Y����l��6O{`@�<^�w�M�2�MR�$�@m ���~���2��r�pS���Q�Q7���d]΢���Uk?xd����ҕs)>6������d�_��~_���u����G����Zsw��:�����������H����§��r洝=wƎ���l�G����}�u+�{���C/�;�p�C?j3o�\^�
�RΑ>^H/�<�
�T������3�95;i��ۧkOm��3����킆�u+tl��c]��A��ze���bk�בs���e��-k���M�x��
��N�w��E���GU�:}�^�����]�>��g����U�?*�A����Ս����v��1�o؅p�p�|=���I��ϑ4���6��x��g��-�={�����rF�~R�Y'\sd��������G�h��!7�	�����ٺ�ز�c�y�FG�C���U����p�bP��8�_a��]*��?�EY�<:�h�Cx�"����`AwC�������^6�����J��SF�O�p ��u�Q�DV���#*��7h��n��I��b��L�$�s�� �rz�9���9Q,2����*�~6��Z<R���o�է���7���g���Mۺ�vWہ��Q�+g�j���6�8o�޾/�E�*�V���1�T�d` e }U]g���r���Q��)�)/̏����.�������^!���Q�l��g_���?���3����̔tؿ�*'��b���v3��d˗.�ʕk6w���^8k��i�ِ��cU��׵Ɣku�.-Z}R����u�W�������)k/�D/�*��+�G�͐z��v��|P�N�k��[��$�#6�e��8;� �~����ܳ���L�Z[�@���7^����}[�pIΒ�J�gGr��r�*��V�Y�۵�ښ�66�`mӺ;�j'�v�%��-���6�q�k=~$�m�V�"�Y�דc�lO��O���⛫��*NH��9ژb!��ѿ��13�t�qPT����&n�+m�̊=z�О����j���y[d����Q����NF��,�����]_G8���C��LL��t�"֖s(ٻ,ޟ]����o�ڏ>���;l4lX���luO4zr��r�ԛj�����p��V���ܴ�x�H{ᆐ7�ua]	@�V�˲��������%��T�s����둵�qC�^���8x9�A�'�Ǉ'��h�4|��<�X�MO��#���x��1�@�1 ��8
|�R�A[7^8` 8'��5�tf'��P�2Gޢ���a0��B��Gʎ��S���L�7��hp�] [�f��LY8N@��XVbuJ�"�p^
�O<�QV���p�(B�8���1�Ư8�}`\.�@/�-G^ħlr��i2��BA�ϴxM1�Q6�yT-�l[;���[������Y�C��Gkv�p뱜��]k(�t�a�����#��;f�.Zb����B)xK=<_�����p�*G�p�^�U�����ExSZY�䄙�ᝇ�������7��ذ�v���lna��u��P;�����uڻ�����5b�AO��U:��>�F[Ω�~[�]�i��j+�$G�����%O���^'�#�h�xN�9G�74`��������UgfF���YKfn�u�7�����ɪ�58��m�>�d�|�.���M�}���t�P�Z�e;���ڶ��cF��\�'�x�*��~Օ�9�o����-�Z�/}w{rpkM[Y�3&'޿>�cG�j\&��m%�De�q=�:mF�5ō��3J�mNȡ��CH'>Ύ#���`��|�ϫ�tpس]9�{��]��봎�V;�H^��ۑ#�W~y���&����)��R��ʍˡ��̴-�������w��X�1i��D_|c�d��$�v{(IzƉ�K%�@7���BW�De�Um�%��ۥꟛ0 l�!c������B������{\����8�!/��(�_L�]h��o�'����4hv3fG���}��S�2<#�7���x:����3Gs���Ѕ�w$Q�j�(+c�G^��0�n��+���Pd���yM��3L1pE~���|q��zܠ� yB��|�Ð�X���y
َ���_�,���8x��J��F6P�,��8���Ex8tH�Jqc������H�>��C��#y�m��Cۑ�2\���?U"C���_�A���[��V;�ّ�0Q�u醟B�p�������d2�8dDV��C�8'��B��x]�TN�X��ڗN�1�h�~�̂i ���kݻc����1ʑb⫢A���Ԩsh��-���/>���ܲ���-��6�ݱ�;�m��m;�ٳ�վF�#9i��9��6�~Wc�A�c�P��������t �R�!���Q]�\[@��]�\�>"�(�kU΍c����Cz��-������{���63��ܔ�?�bs+K^������l㛯m��C������Z���d�{=kJ8��c�V6+�!��)�(ZX�@:���̼�,,�Q

|Ig�ͷAA��a��D�"�x¡����B7�������y��G�?#�Q;����S���3v�4ķԆx[�����yި�Oe��R�8`au�����:KEHG�;m�z�����G6u�e9d�6(q�(���w&��{v�o�g�T�rQ��ϻ�EK �,1��"{���w��Y�!��䍧/�@q���v�6���αMb�1$���H?u�m@|�a���ξ%ϯ�s��8a��@#oȄgff�c�#;N��l���j�1�ޘ!�N�eey��!�:��_J�	h�ٹɛ�;&�d����e�W��'.�wǐ�:cx8�H�,���CB^�4�'} ��<����uc�����?�9"�r���A^�>�#R�̛q!C��1'5❺��b`s})��h���d�q�*m9[��o���Xk�EEi]\�xsn`]T��)k4'�o�UP�V��^Wf]�~�{A��!�|䄲.'O���E�+���8�C^��8=�f��}��^���n���m��ڎvwmR��4�m�؎�ϝ;k�r��6����ك_��ֿ���=�֓Uߎ`��C�|x���<�ý};����اWlay�z�q<f�g��^O���7�����*���s�	.�yu���+�H���5�'�C;B�rr�	�����A��`ڍ[r6��Z����N�=�K�j=9�;س�7����0:6Ѩ�ai��K6�����(�����r��Krl{r(�$�mhqю�uq�,��]8a�$��{}r�N^8��0�� �3��N����<�c��Hm\^�do���s�K�팜2f���v�Y<bJ
S�W�2��L�D,f��e�7��{�)}UΝ���޶�����g�X�R�7w�r�gԦ+�1��F�����V�-�cS��fK���6Ay���آ��Y'̛�,%8^���]���!7�ǖG蓏s�18q�c������h�^�E����������	�w���B�;>-���tD�C�S�8x'+:ַu���>�_��V8C~��_���C&��4�x�����%F%����(.��e��y��gd����7��M�����&�Č�8]�=��Z��'�	pb�,u<$��@�Xn:%�y�Fƥa�A�W�t\|d�,X�8�^w��<2��]:�Vr�<%����ֶ7��ޖ�T>Yf_+Š����=;�`�m rjN��M�N >�iF|"G�N
���(��*t0��pl9BO8�����Jj_<z͙0��I����[_�ރ��y�U��43:����[�|�3SV�o��;���7��ز���6l��c�y��g��[>���F�L7��V���=|hw��F�����5���K����BR�V�9S�ﳊ�7ڃ�8�7 �.y�'p�����"���^}搷^�D`UE�P���ꪕwv�(�'z������!��V���V��)<����5�t���h���[��oؠӵv��`^��E��#q��6�e��-5�v]1��gqV儨�|i��ٟ�]B1�v��HD��<�}p�򏟣��ڑ�
�(^i'�c��:A�=t,=�d?y两�~V��u����w�j�Q���~[����3�����K�ls҆9�g�}�.}���x���u��X��������[���?�k�KKގ�]�I�T$�v���V�@,�HY���������1!���SsA~�4�cm�7!9�!ˊr~3�}he����q'�'��h�9���i�tD�.�x1w.dt�x��K�pc�#�C�#��Rt X��Y��CX:�I��u��<����| �|�"��+x��tF �]v�?f�2 ���3a�B�_o128���r�� D��&_��)��o8m���F^=�׉7�q�yD�S�ͪ*0��E�sg6���J=�(�e��ѐæ�Ӎ��]����������ǒ�$g䐁ں������a6)e�7&�i���4P��fp�R'�+G��^iW��:.�\�H�B����� �!����]o(���*̚�������������;�ځ�� ����kͳ��<ٴ)�E��M<]���X|���&�&]�]�m�7�{����ܜMOM���G��l�V�=Ty{�V�f�dL6|pw=�&2���e�ЧBƼF�8G$��A"�!��Vg>u��U0�bѦ���+�`��Sw2�ɂf�T�Ou�>���u���:�kB���������?sFt����6��1d=��'�� p�y�ͦ��2N{����v�l���[���w�	�M��_�䳪"���t�E��������IB���a��]��(��^�oIg��Yg���?[��w���o��w��W��/t$g_$f���x��q��������W{��u�%�Ͼ��]��v��)+��-��H죟~l������/lo��u�w��ma~Ym��ކ&�a��N�A�Et(��~1�6���~���Z���n�qs)l��������a���R�c�@\�4�t���5!i|[�����	��l�4���`��_���N�`h��d���B��돍
���28�ÞJ��KPd�8�Hǅ��e\�z0�c:E@���q�rF^ܙ�&�A��4�����$w��2�gp9QJc�(p�J�!���	�1H��xQF��U��~���1Ji���Y���x��6�<���Y4=�A����pը�)9aM�kX���^�ko�ju����g�Y߶	��{�È��s�6��bG�� ������^���6w��M�^�1���G�Ģ>RFO��������>;�A����2÷��=����ړӦ���L��w޴So�n�gV���9-�s:�k�l��7֐��A����w���(��o��*U�c���n�J�*GޑO���T�f50W�u�lP�ٓ3���y���}���U�;�6pR���GzRX����q0u���	5�wz=;P�`W�9h��ٱ6��5 ϔ�6-)��HN�X�ݓ#>��h��߳�x9����۷9l�0�Ma�؂)&�$�dvޔO|�˩-I+o�a/_�ʢl��/�cv��cs�fa{Uy��уA?�q�~�uࠓ<2�Aho���g�t�5 ݩ��O�\�������_�ӯo�psϚ��Շe9Ern��{��-_�h�����?���w���;r¶�͍Pe��o\�+�g�����p��vl����翰o����/?�çr~ןپ�	9���s���E�1���+�)|��Q��&7�ԁ� ��#�g�Ҟ��6���pW8�SӾ�o`�������l��O�����	�w���8�!x49�����c��0z�wd��0Bt ud��
�[�H*���A��p��B�bhs�Q�L��X&Q�ᜑ�ّ�Hc���`���q@s�.�A��=�E�_E\�+iL�'��D����o�COd ��2��Cq=N��K}A7bYS�����mݹkO��i]���{Z3^�qt$�G�T���g�V���)�s|f�&o���̱w��%scn��Ν�jsR�k�d�y��/>qB�S���l� +��#�����|	��u0,�~6QN�?0h��1K����P��U��.�uM��)�,k����������۶~���=�#�'��W��?Ӗ�R��Ґ�29����&��rΐ�նڑ�*��v8"̄�,-Jo%�,M�-1�G5�B��L#DB��g�c���Y#_�(�>���%��1
��-+��^V$󊜢SK�T�=���0-gX58����$�xl8aȈ�Ԓ�֑��U���G»�A:t����h^<o��]��=��|�&��g����rm!}-j+`"�̰�m ^����ٯt��$��.���*��b�1��k��be�g_7*թ��x0X۴��O���2U�u�ߓ�ݼxƮ}����v�v�s��M[{�����=�//�˒�ʛ�����=��k{���l��O��g?���G���	^������N�^���l��Bfd�:�md�`9ѓKkM^��bvQ��g�ˬ/�M�ǍD�+�.^����F����ϔA�M������'�O���@�uS�:4o�����t���wP��k�w(����|���G�΃����b!-�e��B'g�9�|�sMNgC�".gb0�0I����lA/��8��Ñz�G�:���N#�|��Ϸ��N �a��c��8$��Q������pB��f`{w��W��2��&���j� O��Zcz�gCXp?/�Y����#GK�4���[6�۷#$,F�7q�t�\_X����X����)����Q$|�^X��)t|NH��RΑ���
"�w�1�:�=�x��#��*�кr۶��f�;r��%�J�t�m�Oר��on��o���gC��*�BG-�>e+��XW�֐�A9)C�}�x�h�$\^h�1\[�٫������6`���P0}�h�y!m7�xd���e;#}��Ņ�Һ�Ǒ�����KUe�5O���s��J��z����}woG�U��1��ܾ1��훣Vs�z�w�Ė߰y��OBYgpd���O/�������rÆ*��]���7�s��C>�M�����п�pA=����8��7�X�Wp���o��B���zC.��F�-���[���Y�s9?��@N|�6M���%���/��{�m��7j돞XgON����}�.]�f�����7wl��7�싯|#ے�W�@m������3�U���=���)�ș:�h�I�$Ig�/�� K�6�IG6l:���ΧX ����[��[� gO����ES�A��;A���!���C�~8q��D�Ec�����wP�t��::�?NR�ht�x���°F@�y���EYdC��(-c�A1��-�s�Š�球,���_�#�,��	G3��y
��˼��"L|�Γ#��I'tF�A'��A�����8��Ќ�qH����uF�l	�teS�rLuW����~L�o�@wՓ�V/�ؖ#ɛ_8b����P�6��'�ڣ[�lRz���J����֣Ǿ��7&�[ijҎ��6�;橅y�����o,Bfu��e�C�����1g�99�G�)o�ŉ����6�=��hGJ'M�0�U����wm{�uv7�0:V��t(��k�o�����y��=��+�V�R3����K�·��mK:��ݏ~���TF[B�8�PyX�&mX[e�8T�s+��13'�G�ɡ�V�w��h��i�,�#��B& �0i9�nk�$7�f�Q6kU/qy�NO_c1~}n�jf���wlk{��v��2�-��u���8�������+�~�	������[��l���v�;Z�6����9�l���_o,d�nb����U����'=Q�ΊzO;��d���kW�C�AWd����N�|�!��/�g���xef�����X::��u{���^�����ۼ�����q�ʑ����f��;{����	{�ŗ6X_�SW�}��>$�UGlm�����M�ߵ�l�f����f��n��ie��"w���x}1kO{���j"��z�P�o@��b���܂�)�	���q!u�"�=�����9�?�8a��F����O������bL%x">�~1X�+D|8��<�ț���ˎ�Ctc�1:<��P�A�1
>�+>ҽhS\����|��A�NG Ң��7ydh8:Y6�G����Nx���O��F��SXiί~�O��A����q�8tu�ׁq��=��|�n��V��o�bqy�}`-���'c>��d������-[���T���{�{�i�=�k�v�g���_}�j�����u�--��ٳ��䑜�#ݽ����|<��!s���&~��X�GZ�.ds]�M	�G��y���i��5�!
r�Z��#���U��ViV$��v�>���m�� Uf�������ɗ��ĺ�V��0S④�N��CG�li���o�y�S9�#����v��ȧTg���֗�3��l�/]����.����	 S���;�C� �Y�+Q�b���P��=)4`5��q/�Ø�8�S1o���ڮ�����f�lj�i˧�laeѿP�þ#'��n���#�r��3d]h�'ߏ�2����Ȗ�a���j�s��ƫ����Ȧ^�l}�P�6�YkH&թ�=h���X]e�*�������]�ɞ����B�v<ůUE׺��`�Х;���tf#������,1�>{t��maiΖ��L7�G���a�|����ڧ?��=����ζ�� ����{�j;���h�e���I^|9���U�[9��o����dߵ�^��kG6{�͟;oSS�TM�4}�`lS���#t�c&�G�CQ����jWN�ds�Ξ;��5��A�x\�����!l쨞~������'�I� :m���f?�)��#��S�-F������>���2!�c�F �P��*��"�r�tqv�n�ﶹ�S:�Gz���t�0N�>$	c ��:�ھ�8.EyCdu�µҸ��GC�b���	D<��j�xFaw��()��,s�[�yj��������Ꝼ�}����3�Q������򕫶|�%+�'m��#{x�+{���֕�1/=�7�l��{����葙��6ԝ:�Hsf���̊����v�_�Ŷ�>�@.�=Ӱ��tދ�(ȈAg=zdmY�$xǽ��@�i��u@�?ҍ���8�Hv�:M0CC��'%ę�!����G���h�q�kep�;lN+"<�UZ��A�Q�|7�$y;�e����utfm3}��X0ͺ0N�k�ݮtU�v�μ��M]8g�fS�KO͚��tZ�:jrb���+��ے�r���P�/��A�Ҳ�&M����ڥ?��߳�w�M���� t�ʬ!c}~��.\�Wn؍k�ڍ�/�޳��\��M��/g�o#�o�խ?uߝ�O�:m�����m��g���������/�����#��ڕn�F�~����޺{��ۛ�9\��d]uV��s'�M�"K�T��E���j8 ��P��s��d��g"?}�:����/�0�?��t%�IAJS���o�e�/_��/]�����?��m~��ܿ�:�O6	ȁW��^�֕�58�[��~,縤�����;�>�X����H��{8;is�֗C<{�-��$'y��W!��F�W�� ��S��b_��;O��O�8c/^� G�):q����opC��9�$�����8a&��D�36M���*F�Y1f����5���g������O�jv�����<:�1�C��D:4<b��A"ić��1�Ν�I��P�FA'i��XaL�p7�q �)�#7�.�]�q
9p�0��NTd���Q���V�E��Q<�8�7`�'x����Ne$�[8f��H�L�<U99|�f���䩮�3e�NO��K2�W����oDY�kp�ڲ����5�}��>���a��i6`��]�˖lJlm�����24�j Wh�l��`�#_��<Lȓ3�{�c��\��1=L��چ�&�sD}-�I2*�̓cPe���qr�Zj��!�񉝁dg���)��� h�r���Y
^B���9>o����ԱK�@x{d���d/��{���uh��g�Y
k)oCM�Q<��K��\�A��~��VD�֙v��^�a��u��h�������5],ĮD�����C���)�5Zrx��׿��n��3�[�Huޓs����wE{r�O��K�_:^?������;=e�>|�^���B�c�d�����ˁ<Z��Gv��ٞ}q�z���Mӗ_}��j���ȥ�fM��q}� ��G�(�3@���f�)��aW����N��́.}��p�:���Fc~ƶ��mS���7����}��F�$Ǒ��Ո��T�Cj�U�Y��Sj�la1���oY��GiÉ�����~�N�ęS���v���l��e�����ϰi簏'�������$�*��kaI��]ᦛ� ���x#����E����=�?�8aF0�I0L ���p��}�Q'�E��L����?��"�N���??�F#�v����9�.`�,+i�^�'0��୴�(��=y���#��x����|t�Čsc��ƌO�?�@��������@9k�'�'d���/�t������u6�|q9{�Y�f�g�X�̊�e���6�A��S���#8f�:-ݓ�1*�&��2%2��'e`Hyzmk�.J����)9�3S�6�C�i �;c��[���4�r�2D�#w�FQ����N��?�D��W �:r05-���]@�ll�Z��%�(H��:�P�!��f����a�<�[�qO��)D�]8�����;7m+o��NHm�u�s(���
;>�]�1^x�'L#�;�^��uy�]�H�����Z�9t��	ex8�ɨ��c��M�Z|댘�I��Oh�&�1��_>�4XW^_��v%HS���ۯ۹+��GK6`�ݳ5��S�����ʇ�مWo8�R[.�־�������K���m~����?���]k(}(�S�3?���{���:�U��vI�o���~�K������"��	�R����������g���䃮?����VW���_���]��op�b��yif}������6�4]�Sr������{��x�=�z��Þh�n�.}�;v��l����-��7Z���!y��p��En�sw|֎�<�?�|A�0{��:�����5cp����;�8af�F&;h���S8bud�2��m	�t��t����iɏ�OCp�x�
��41�␱�GX##�icƖ3�X_|Qv�H�H����i<��X�98���1/�@��<�/y�c�v�6���'>ɻ��?י=P@���SC��uvv�/���#6b�u`3|b��i+ի��c��[�}۶=�����xsOw��6��R�|���������
���:�Tx�893ū���7z�:��<dB��̠�B��G�P:v=��B����uE*	��L������bJ���|�5muk�v�{�7�K���i��8��"'L�:M��W���<!����6T�����oMO��;o�տ���]�b}9_��aP��(vC�M]�5btFwx�	�B6Zu'�BFzp�BD����u�8�
z\��(�0 �tì�;�Jf��I�ay~�.�>c{���`k�!�iH����-^y�>����K|��۶͵����mn>������g��;o٥�/����ƞ|���{��_Xym�z���������ၜ�~�7��m��ڬ/"��pU->3��UUu��]�Cg@�qX\��o�ݠ�2<O��3a��>����f�Z�)�c��w��`�����n�b�s��p��]x媭�������AW6������)��&mK:8���c�~�}[~�=�����Ӓu���n#��~���G�s	D?��@�a�����:#'�4l=:�C �����xp����p�`������rW�;I�Ζ�\�p:��(F�9|0%\���PW:��A�0w�q���H�\�1$y\����A7��iy.�'�M8�X��)儬;��9���F�Q���|L�s��q�q���x-Fg f�F�:s��7��cg���X�4ё�G��O��XMNؔހ|�ŗ�0]�wa�54(������p�<F)�=���#�S���Į��JM֭�8��T�K�C
���^��!AnL�����GQ���8O��}�T�Syhr�O�r4�.\�w?������-�,��ܬMN6�%���MqCT���&����Ԡ�w�[壊�����z�����+���[>&i]o|�s�9����T��YC�U+[W�'ګ8j�*�oT��.��F:	�q�u���W8�3�k�f�k�cFN�J����^X3��V$�3���c;l�!^옿~�^��#���k�5��7���{w�`g˷��ˑX8}Zz�l�Z�n~��m޺k[_ߵ��U�ؒò��6Þm��S����J>��cm��x>�G�};����D�Wa�L}��Gꄳ�]o#��5o[��@��-��U�af2�<�?����RW>�&ޑ#���C�?h[W<�6s�]��M{����[��M�ƣ'���ۗ�l���<��{�ڷ�̬]������}[z�m��S�oN���U^�{ �cm�g>Eŵߜ¯�fm/�$P���c�9X���O3��N~H��}��}��	�3�40�a�t(:$>�������k:_|<��?G���k���)�}&Ae���A�́AI�+�(#��#��1,�j�v���rbM�^����Ȩ(/�HW���#J
ZN_~��Ү3�s�<Sy�˲��(��?�QZƏǅ"O@���5Y��wՑ~J�O�쯮�p�e͡x���߲}��kk����7m����5��^�XC�Ȓ��+׮zؗC�V*�����H�O��i����Þ\09���V�6�@?�w����,j�������8h�,=��1ۃ�Ɲ��=aA�{J����Bٗ,|J��ٳv^�P�Wk}�* B�)�GE�r �ĆtrZ�AE��^vV�WuR�p�.��w�ʇXcqI>��/��gW��C��}���Y��q��fM9�����¿�-�3�Ո�.�yD�+%xG�+�e�x��9ɶ�k<�l�Z!Ѡ~x|�L/1t�������շ�/�l/}�{vM�Q��{^mܹm�gkj�C9w�jպ���z�=�s���?��ξ�uԘE�rX��VY�)��S2��Z;�X�S?�j_ͥ%[����kB7}_,W2�(��+"/q.'�!d���l#�x���ٮ�AMѮ��OՉ�*���^YZt[��>��:>{�]~�M{��~d7~��5fl��C�/Gt��;v����,����*;��3f�WV��h/��_�̫�X_pO������ܭ�xb+x�F{}R���v�V��ڼ� ���<M`#Vց�����$�����~��4N��'N؟dG��bx��s1s�a�n�;)��VZv�<{GT>�&N�?JQ\:�m֦���tK�Ǒʜ�u������I8�1;��f�0
��\]cl���s#��px�Ù���B
H��!.�b�3�����L�Q|�J�3 o�
~���z?��ϐ����i4s0�i	�
s��HM6d�{}�m����-�:*��d9���ll���Ƕ���U�]_�s$#�kp����#��mnn��
G�x�l�韥�W�Z_:�f@\����S6���gޥ'�B/!Z��r)B�p���É�v���Fۢ��C7�EH8�}�y�pX���<^u'[��U�s`[r"�������Xu�eu9,Bo{֭OXG͢+gaN:���k��rR&lw�%Tlg0�����G��:�Ϟ�Sհ���Ξ=�����?��=���l��olb��iצ'mae�&����=8D.���q�Q<zr]�w�ŕ�L��:�I��C��ä��^�p�SF�3�6�A{zq�?�^���+o�i/����YZ�g�n��O?���Slo_U���q��������u��dE}�5p�j[��(�a+�"�C�֩x�0����=�é����rJ��~Rv���/�C�1�um#�su�_��ǅ�8�i#>;��ӧ�-�x��3�\�֩nj3e֋�J]6r��)�?'g����᏾o�_���坏a����ڷ�m�͊��PNSGz?�]A��Y���i��C�y�����w��naҧx=<R_�c�b�oHb�CR��!�.t��6��N������D�7����s@+ʏǢ�/�O��&T�Es8�?wȪ�3��{�lCw�� �4����c�����x)��Jң���E ���8[ܥ�6ō���(��.^֝ wt��ƀoP�ؔ�Єf�H7p�C;S��/����w�:ȃ�Ę!�����0J�����6�l �)"Fƞ+��H�C�q��ǝ0�	�%n;IZ�jP�]�������b�;���ߝN�ʄ����Ls�בIw�ϫ�,o�����^B[�=���ڄ(逵`�MJMNt�\�V���U��_����v�7����<"7"Ǻ/�)5�$��� �Hw!s�M��?i{��H?�e�t�d�;��%��h�� �q�T�=9�_|i���O����mrCEWN]�f�����	���-�>mo��5�t=�枭�{h�rb����K�읿��]��V=�l뻻���f���m߹k��ܔ3��6ģ��5����ik^�.�[>w�r\��E����3&M�mj�#�@.d�6:������#�O1��fU9\��J~���)ʪk�e9�3̫}����S�Uڇr�>��?����o�hs�*��oq�~�bzU���\_uu�z���x+���2�ؤ�*�~ԗ�ϖ��Nٮ��f�^�o�Ֆ�y��]��;�����A_���ǆgʏs�l��9�q���V�c\��HCo�-t(��w��.�<i]lB�������7��ZC.��4��d���ܶ�?�G[��Sۿs���p�s�Kٜ���h.\�l/}�C;���l��9kת�Qs��x4�r���{�6=�n��҆lq3��p�$}�����b�L�a�����7�7���x��p2��@q��Ǣ}��y4�N�ħ���r >@��D^f)G�0lA1�?�:�	"B7�:�<0��� �p��/�-z�G�\c���=
(;��뗋x)��<��x~����FAȝ��iH�����X"�=�t �SR@��Fi���y��âs�A�i(��6l����f�ց�Vor�4�K9�dv�g�t��b�֭�>�wJW]�F�ן����uR*��떜����vI�E���%�jTtE� � ���x���D�:By���I�))p�Q�c���@��= �U�(��P0n�Кǋ�CʱgF��x͎䬲辥a��P\���l�����������l��S��ܱ���9��}�;v���݉�Z&'�{����翰u�K�[��ʑՠ]W�����u$S�g<�)��[��s�D�G߾��e��GG�ˁ�I@ ��"u��zm���m�Wb�J�I�쎿��Wv��_�����zf2V�^�}���Ӻ�a9�l��M�u�+���
�����(�7ǚ�����]���څ�ޱ�+W�H4{rt�/}�m�MK׌��6�?���8j!g�)�9Dx\'N��@�4�|�[�WLI�/g� ƍ���Qo�c&q����z��Y��3[�^*js�xh�H�ִ�a/��GvVr�^���nb�`��	o��7'�i���w@�;l�.q� ��.��"���~�nܰ2�G�y��y�w�&y�}��Q:�?8q�������k:"k������u�s��t:&����` �����J�E��8 z�_�C>���o�!��C�'E��q����
z�9>X.@:<&.N
�}�.X�Y���N�w9�x��*GGĂ�D8�����pGS4�		�ND��1v��H�:ҝ^A ��r�:@��f�&je���؞l��~{ߺ��;U9�yaI��b�#v�G_�@�&4�2{��W�fq���cO,��ϝ����;�q���3B�UV�5o��9X�N��Yr��jPa�S����Ы�q����|`Jg��傒}V��Gf7��Zcaz�Vff}6vkw׶�Cm�a9�_��|�];�r��}��=�����;����r���+�x���۝/?��_|a��n���{�y�Ԭ�aW���r����w�>�^�T�����e����5@=�5n@����G�� r҆ә@^�k�_���J�h7�S�RgT�eY��,�2�S
5�D��j�A�֑#���?�'�[{l3R&��� CWm��v�g}��ͦ��l�6�����U�����U�P��j֗#��R�SM��t�V��^��Z��24&%k�����ao�O�z���B&䋶mJ�.���p�o���s�#�>t�G#���l[�$]�>���=����Ć�ڔ�yS���n��l�/��l��u{U2.���UO-IΚ�iaE���Xs�+��g��Q�ش��a��.scK[Ff������) �����x����?�{8q���c4ȍ<3b<�dsלm�;�0t1X�:)7^pw��P0�XJq.a�h�����7(1*i��b��+|��0p�;�d���s��E>]�p(����8�bH����qcV��?�((�yT���4.0���a�r���v�z�ᮽR�
>��;�tw=�"�/g��ųƺ��֞��m�`��$Y��[q��đ��"�&Ѝx8.h���}�(��h���-��]���6y���E=ș���U�c�YbfB�0��ZȞ2��Aᡣ���t�3���v���p��kd��Qw�ߗπ�l**���j`������S֡�4�V����7^���{�?n���#{��W��豵֟I/��i�aIQ�}�jOo߲������j��-+w:�@NU�Z�ʤ/�F�Ǐ-�*8�=�:������9wR�Σ���V�0�*����(qb�=���c�N��C)�Z8>�o���}�W��o��n����͈ ۠��F�k�z��.\:k��zŮ�|͎Z=�����F��<��ObRʺ��`y��~����_~`W����O��}����se�%�Ҁ�:��_a�9��"ڮ�?�		�OG�h?#��$�xp���B��I��BU�ꕢ�쐴�z��|��$�8��֎�ZOX�W��ɫ�}��q��sS֒�J�cV9�+ .U6�z�ŕ]c��o����	D�cg�$�<��K�pD��� ���'3`�p����a�pt�#__����aQb���P:g �c���P�tl]�~�P�8D��9��F�7��=�R���KF�|s����4 �Q�7���è��(�y=�/x�}��㼂Z��"\�@�3����2
�1W09�㚱rH#g��I,���_g�4�XiG����K� �9?cg/]�˗/��bmk|����օ�G~rnط�;s7�8;�S����%�mNZ��}����r4;+���y|�El��o�v�2M���}!��<�FB��L���������Q����3���q�P�,��5uΌ32��G�����ı�EerҌ��y;��x�-9�u�^]�'7o���6�ݵ`�#Z����ֆ��^Ϛ�u
�T���\�>,�����tO<��@��rf�K6s]��苷U޶�Y�v���Ü�����W���4����e8`8�x��6�#���,5�{�.�lo���֭�_8�T�r攝y�U��z�^z�e���%+���_޶����P�vg^XW�#gw��e�*����|��^�f��Y������U6m[q�&��x?�]*ɲ��:�y�8�=
=D;�p
Ү�_��6���p���Q/���ʊ�4��^K�9��ئ��V�el�kTm�������Y9a3�\��줵� �u����}K��ri�| ݻVȊh��}H��G��efWї��u�� �g����:�;8q����#�%�����~f����M��is��N�A�� ���N�t:J�10=fh�������A�k0###���$fJ� ��q��p�(���= ����,D�ΛE��-��@&'�~�3G֨4c�ҁ�bh�}��{exuf6����z��C��r��x�T�	��������CN�_
hc��%f5`�k��i�H���#���v�k6��]]<m��k�:�� Ϯ�ʣ���%�`0Q����r/}ԫM�"�)�Pi�*�&�n��W���7l��i�� -T{V�}f;woك���V?�܎�5�Nӳ6!]�(�C�k��Y�D�ñc���0��웻*�^=���z�N�3�D����a��3,���ɕk.���S��V���m�/���Zo�u�6�u�FV�1�>�d���*��yerFuQW� �H·�F��rC�3�=���f���m��5������l=��q��0x������t��ᐗt��J<m|�Q9������ŹC�Oq�&x�ݘ���{jS�i�٥w߷����f���m�ִ�ږtv����ml���ǆtQ홵�=���e[��{v��߳�?�K�R�<j�]N��A�FW���_�f�&׏���7�MC���
3�Ѷ��t�sN�n� �G)G8>ˌ>Ƞ��m���rёlNIm��*v󳇏������g7~��v��wm��%9�MYfp�1E���::>��=^�Ꮧ�x��������kT�;č��$ও��s�X��<Ș�bҦg:����m�N�OdC_���O9 pf���U�-J��y\9���'Lg'`�g	�n~�Fa,��D jr��DX�6zDI����C8֐q��9�2y��B�Lt�C��OKǬVWyJ�1���GJ��@s ï�}��a%萌~��?��|8u�]ъ�^��e��:	���=?�;C���U�5��H��7���?���wm�Z;��b�E�2i����x�6���%��(m��}�C:���d�.��]��m��ګ֘������ڵ����ߵ���m�٦oo1sႝy�-[�1y��iA��Ǳf�u�E r� �1Ym�Ȭx֒���@��uD�]���<���R�Ի;>{�V�ڲՏjOt=}j��e�a_�r#Q�y]��x�lnvA��"|qn�͞7ꇅ�}���Å�v�;إ�~d��/�|c�!��:v~D�rF'���i4K�U� � �9G�H&�~�g��;7*;qR��������v��v�mB���/ع�%۸{�>���n��U9�l�Z��ڠ;��߶.78gOIn9`�cׯ�pfڎԟX�<2��K����#�]9axR^O.�9�R�C�xoS��>D^��v���N<5�\�ǶH�U]�؝�n��~fo��_�u�LOۮ�"[���t�3��(�I=��͛�}��M}s3k���BO�_+�����!�R?�����HO�����&�8a�	!&�8,p�۷o��,�'7{���,Nѹ40����@3D�h��;���'7��&��&?��H��&�؀���k����^:�Z���`'S$J2�*�|U��n������Qoj1`V����j����5�����?��r����	ęP�o��N��pu=�) ����#60N�o�0w�86��?�-~�������5���g���`���6�xf�֞��7�:��u�vy�����l�i�c{w�����O���Yk^<m�~�.������[g�e����΃U�z���W����甼��S���6���v������<�	�1�*\��6�C�"�-A��}P�C���dO�"��� �^�2�h4�=;�}�������>��*��m
�Q��'�_�Áoϕ����vvf��<��M�3�qyc��!'�O�l�۶Ө��Wn؛?���~�u���X�)��夹#-���%��m�D7ďd��9��3����x!{A�g�
}��0WRR����|/Rzj����q|�O���~i[_ܴҳ-;�Mٰ�~/Z��tU�������v�/�k��z�g���ܜМǰ�F����e���3ھG�5��%�Cޔ1���?A7u�%<*/��3�N�����Sm�g�_<PT�c�<��%'�·Ue'�I�ۣ�/#Y(/�j��=��&8�G*<�S�̙�>V�G��V���aTn���[ƍC���t��q�B���(d���bA(N�(1jih��|��A	G�x��/ފ}�è��L#����H�6�K�"c����]�lޚ$<-C�#��:a|��ǝ�`���T�o�����b6!�`���߱I���3���Z�/w<��c�:d�+���3q��T�z<r
�A�xf�8��<�d�[;۾���AW$5003?m3��G�C{��W���ek����ڪ���d�\��+o�b�\��8�g������m���b�'���zK������y#>�r�i[_2N��Z�Y��RD�!�뀐�9SI��x�_��x^W�h@�K\�ޮt���u� zk�=��ƶ�oy:;}��So�i�S�ּpƖn\�7�z[�V�������N���l[�F�G̚�}��k6����_��^��}�X\�]�B��`Pk�v�;��G}$D�\g�q9�WďdB���q1`{���G�E��F_X�^��$⥆o�|�����m{_خu�-�?O�gvh��no���f�>x�ϛ:�ړ�H�#���@<_G���n\������C6��@�'��~>���G[ 5p�O���#�3�*W1_�C]�M#[�MH6�_�o�I&n���B�>
�Q}RX����ǊN����.����K�+�4�e�>��N^R����ş���8a�	�N�vd,�cⴰh�u(�A�N|X6��x'�x%�ŵ�F�g��@`����00�D��_�">L5�tU���(3�n������B1Cg >����7��F���u!gM�oS�+���q4X��]$��b�#̿�� �H��^�?t�2���',�᛼n����c�'Nfgg��ʢ���\�m���Jϵ�9��r�^{�];w�=�{�n~��y��[W��y����Sv��)�����/o���w�u������\7u�[�#[�v|�~Wu�7�o�Ӡ1��������笫G<0r���܄��V�F��r����ADVf1N���Ҥ9U��{r��;հ�Ҭ�^�lW?x�^�#���b�r�n~��={�D��2��0�j���C9��o�f�����;o[�Ѱ����;�|�0���Ő�R\e��.�6�|�(��O�FZ�Gf]#w�N(�C9s���ς}f,����?N��mS�߽��ZwYIN؄�v�c76'�LOکw߲��WvFr�VV�����pH�uf��Ǽ/!W�M�o@��B�@G� ��k������C�4/i@3������E���l�0�XjO܏�R���K���>=IY�^�0q�e�� ~̦�H�2y��[c'���"�B���Ӄ/�a ߱×�~S�	����v�1�;<��Y16yŉa�W���qr8�a�N����G{2��`]�H��6��_ |�'���?7dn$q�0JyCÀ����S^9|v@	��(�yԙǖ�Y�SeІG𔆑����d6u�HB��#����l@�Ȉ�,/[�!r�@��QƁsS��u�����kV�����=9�ͺ-]<o���v��K�����_~f;��]�1`Y]�54Pvw��/��|��m��ذӖ�%K�h_�uY-Η)�D2�́ݮX9��+�lfv^,I3^.��C��Y�NX�P�Ã^��+ �U�Ahq~�C<���tBu�數<j�c�w`�ɚM]9oW>z��������S��ײ]9 ���=��P��G��]U���gO۹߳����fn\����T�!<�)�1�T,9i5�'�a��^c�-t�I�+�8r�9�8�y���KV_��e��-���}�W��ɇnq�ʇ�#�.*���mF�y�ɺh��.v�oma�.~�{���Ɩ�y��� �'x�>��^��Fc�e��^<Ï���Qȶ��QQ���cF;�h' �f�(��[��3y �x~ښ�Џ���e&,$���ȣ�>��Y�:�샳��E9�霼Q��eg>�0�:���� ٦%���}�� :/��t�N��N�����b'θ�3����S��l��3��Cg�� ��J�/�a�q�Sጅ��A9�P���
w��&��̆�wc���b�>x�q�J*�����A�A�|
�o&�acM�����1P�N���x����}&%�=��Ǭ
`�ݘ*�uA�C�TV:�	1��$2!��¸d��f;��/k�|P{��&�6�~���Y9	o������?bz��m�:VV֖�1�r��r�w[6�`�y�c���PbptES�I4�"�0۳/�~�am�r�/����E�[��r���㺈+�^�U臁��g ��"爖N
ڙ�^Т=�R���g~td�M��i��^��g�|��M7����={��-����u6��P�I7,�g�Ӟ����=�������{o��k�YY�K�rj�#�P�g0aֿ0����8_��0y�p�| .��i?ąÚz�a �g����ϙr��#��)/�ի�yr ��f����z�_�rɞ>[���밞�ݱ��g�����$�u��e;��+���jj�.����m@�f�d�#�0��-�>gf��GȊ��:/�I�QF�	 ��NP�I�;����6(�GI$ӵ�y3	i�����ʠ�zۓ��1���'��	�g�}�R�~�֓�O�>�K?b�P�D������`<|�&|�����&�,�?�c����q|g��ݻ����f�=�!G�v(�c�q���I�À��7�x�?^W��q�'��3?�t�Ab]te|`¸�ȑM>qHbz?�ahé�q��b�>(�[�^�u�χ��X��i��C1�bF�}�ʍ�/xg�I>��<�!��8�qkN�
���x^�il1��&����8��љ���1H���O��^[΂�N���;6%�N�����ӏ���~n�W]�:�H�k]p��A����l��V��p̂��T�4h�%k�9i��m魷m�����+V_��æ2�r̨ne'��G���}`M�@�Q>[b�S(�":>��uO(��O�RO��N���t+ɡ���u�ۓ�Z{�$�k��ck��ܞ~����{l���u[�Ǝ鵚�j�:R��㙷^�s�&y'5`Zc�z���\ԧϪ��q�^U���d�)���NP�פ���l�)�8@�4��t�שG�%�C��(�ߺ*-���N�Vc�v�?���?�ľ����|�f7>|��~��-_�l��9q�ڤM�'}���ʤ�&ԟ�Qo<��<�C��Љ�	�����"����v��H'��.��aJ�;~���}��r Q/X��&���A��gt��Vo�r���CWa���pc�q�Q:ogs���{�>sZq�O�8p�A�_���t��ߔ��4��	;�c�uM��M�pmm�ߠ��ڶ�����ucÞ8X�x���%c�|n�5 ��8�+�7��I�*Wٹ[v�	��b��m~�Sy1���0�a�1���qWH�;S�o�wX���x6���rGNNϪ��F����!C�<��6��ծ١���'����t���0�
�xρ!t�A�����I�u��>���DF���t�m3Wgd�VlF�'����������y��z�{r,į�j�뛺2�&��Zզ��l(G��e�_8�����Ҫk�-T�-�\;w�ο��]��C�j �M�Ĥt!�J�Q����H�J��5B^��)��D� Yǉ��|�'gtH��vm[��۲�������o�g���_��O>��{���ٷV�����΄��)[|�5{����&Y���P�5|�,f����:���^Ń;R.�3�z�z�GE�pܸ���ɛN֋y�	S��4�C����ċxѦ9���'m	�,Ml��#{B�~�Ȯ�=g^�f�����.e��~t]6m��{�A�eR� �L�\?y$ދ��)���ö�qw�bF�cD[x������Ƈ��N���}?fI�8bC���Ʀ�����(�4M�������T�A���2�oA�L��JY~��{��
~[��ӄ'�~#�<�(��a��ܱ��k��ڱ���`��8���U.u&?��h�y�	cC�#6g��XMw�1c 0[3b��f�1���\`T��%���kd��Ŏ4��eC�e��5������#���v�.���/��_� ��kt���Y��v'�K*Ҝ?񮁏3�&B��?DFh���C�xL���� !�B&׎طJe����p{��>��=��m�˯���oU��c ;�I�~��ZÞ�f�lye٦M����n���?���k�`a{�|d[��u�u��t�.����~�-[�v��M�(����˪��] �N�1�AQ���u!�8pM�F>���c��.�����8�p�L�*X��ȩU��iI���l��[��g���?��[��?�~C�'��$WmpO��k����W�����lhY�o||9(�g�7fcb6�©#�B̦$�_�A�O�ħ�|���^ f۸�>�����z�8�zҡ�^U��-�]�Ֆ�J�����v���#n��f�����&gD�ȷp����&������9��py�V��u�<#�F]�ܜ������r���;뀲B��?y�˺��o
�-f��2?����=�PQd�����
�SXޞ���y�{����
q������x�����nx�5�� �%!���o�ț�	�y�ɚ����%�-����ma~��|d��ç@|0���ύ�w>0tn\�F�SO.)��[?�{�r���ŻGʀ/�a��Q�o�J6ٔ��|�K��;���r�pxt�j�G���'���'�[���g������X�EF�ˉb5��1�#�M���5�����H�o��x�bp�LJe�����OƞuI>3�:�����}��z�;���X�{$>�9�S-Ymi�.ɱ�t����/��Ξ��������7�D�x1�-:��-�r�^��w��Gߵ�smPo�S*.�S8҂;ީ ��P#"d-�:
�ۯF�JA+�1ە8�^UאdFq�/��M�7��V�W�H�}�����lnI��8�����a�������]{���w�A��䔜��40�WT�+�C�i�v@9΅jI?����=U'��6�#��L���e���4��q�G���c���ř>�f�U�F/Vw}�UmhF7R��5���ToX���t&�<R����p'�P�u��Ɣ)G�� 2�F�x�^7�x"�~ċ�@�����E�;���\�G�������2�L��:�6�!O&��<:�9脬`q'� ����N�"H�mkd�`�+�2�>�+#*d�����yB�ȗ�o�;�?/8q�N���>n(0��SM;�r������	n���L�$w�p�C� L�/H�ﺯ|��D���x�ƍ�8t���p�DEi#p8�x���9��ǰ�'jj�j� Ol���ͯm���6}г!��˱d_�R�nU9reR�@��RYh�����6ǆ���^�".����0��e���	S؝o��W�̣Y��pٕ&?��\���*r�����ؗsՑc�[|��i��ƫ�?��]������ٓ��lgm�y�� :����+f�6�5/��w�����޳ک3֯O����%7#<�^��CF��sYr6S�t��JG$f��
�Ѕt���h1��W�Ex��C�p|���>��z-���y���v������b��͏l��E�H�	>��u��үZZ8V����������ЂP�S:�p���l�
��	r&-D汣�-}g�g��p0F�a��Z.�T��Wq����z��M�x�hN��F��2�&!]��r�P��Ny<ɧ��q�%	�I�z;��{=��������;�hE2z( �PY��0�#g���p
4��򼿉�	��C!&/l�PϪ�?l�4��a�^D��5�E�������Kgf����;`�3�O��Ѩ>�!�_�����L߆{>pℝ�o����V��π077+gl�:�ۑC��߄����g1�(.������M�<dTe�E��1���\eiP���A��|#�&�"��Ĩ�]��9V��!I����1]�3!�;{{����HV[-k*E�܎4��q�&��#���k�b�Md?����]a����	a�E)��}GW>x*���z>��o�E�~�#u� �X�V�����|��X�\���gm��9;���������4���ǟ��O����O���Ã���*��ĎHnMM٩�߱w������޲�̌�r�pDT���h_�	���)�Rn�]�(����#��c0�g�>b�������$��A/���5�!�x���{y��n�HW��!=��X�԰�������v��w�ha�7(�Ѝ��)=�+�hk���"0�h�S:�s>2��?d��"�0�;-�9Ɓ>n��Lp4ɓ�5�8�w��"���nT_�-pX,�p��WQ״Eʬ��*W�p�8W�8~4.�]2m���Q����t�d�ExįB^�������72`(�<���;�R$�:!���ýC����N�P��q�4�&�o�<F9�Z��é��
��	o� ��:�-�S�3��uܡM�&uye��.�.���]� �#�8 �ύ)u�=H]��9�?_8q�N�_�X�0�`3��v�lO�w��JՍ�N0"�:N���4x�}I���4�y�ߩ�N=����c�}��Q�3�;�0��la��[tJ ���~���=�J��k�r��&ޡx;��7y�-,-�#'�Q�#���!o0�K� ���kt�30����p�+�c�M�����EՎ�����U�e���k���cW_}�.�|���������|l;;��>��c_���w��v������;u�M���I=x���î�j,�K��:ς<'�,>0��;%O�@/ '�ş;���4��9ʈr��z��q��We��\���������ss����i��)�	ם���V��MmP���ʂ���5Q@�T:�)G���u����Q��qQ���L��<#���
�Ͳ<��Ҩ������1y�(�e�dQ<�q�Yf�d8 �v�N<�>R)_�R� 9z�6Jѯ(�8�_����G�L~ȕ�_;]�u��<���I_�2�w��_8W��34���7���B�����}p�Fe����Y����O�?�,�?�?��`0BPn�w��]���Mozf���7j^49f����y�������z~W̠���##�-��U:F09� )샯�����@��s��r��	�׫�����ڪ��������?����{k�T�pe�f'mp�5o�l7�ذ=�'��r,U�@�4����C\�b���&�8/�u��ڝ��O���EO�8�V�)�����5Y�_R���e�ӵ�V�&���p������mܼ-G�2|p����էgl�ױ����o�n/��/���k�'�m�Yn4U��T�<�C��y4�i8a	/�OӑL'�8n�C�<<���D��ʓj�+�C�0;����֭���Ξ;=��J�o��1����劳�{�-� �S=fo�#�=E�� ?�u�u>N�3x��9G��9�Bn�7ҡ��)1�B���t���a��t�/oп"�t��Q��;��:Dւ�P�~ٿ���2�p�@�<�N��YsM?�Y��	��c2g�� ����ޕ.����{��1�����y���3��vy�od&�?���q��nbԞff��⅋�[n ���=�</E9��{����a�O�?�8a'�f��#��4#,����ޞݺu�vwv�є�Uؐ0��>ŏ�a�mK61dƋ�;���;�������Y4�a��X.�lW���H�.o_*��=��m��������ғ5�X3���*fm���mί��+6�8��w$#�,��̚�/�э�����+�#������9P`�y��F^�f���������3�rHy��c���w�������W���N\Պ��).7'�HNG_Nj�Ԣ]|�m����V=���m�|��!��qem�>���5�Q�G�c��q�O������O�^�#hPW>s�\Ʈ"�
�,��Z�Be�����l�݆o���.��4�7|��h�b}ᵏүj�dӍ ��Nq �#��eć��	�k��D4��L�f%7t�ڳ�Fΐ��v�����hҢ�D^� wp�4����!�NЂ�,�g��r��(#�8�	�:5�8P^ߢ��Y��N83�3�<�c��1δ����pH���~�R!7��mH����	���[�J���=���r=*LY��g�~|�����--.��>��ጓ5�'t�� ���e�o�?�?o��8��0V�Ҩ a(�Ǆ���{���^�;M> ����#o։��#U�$�i�x�M�Pˁ�����cN6|7i�A��YsF�ܨ�t�{�#*��{49i}9]���ug&�5l��Y�����G�՗���ƕǩ�X�!9*s40�@]ބ�O�<��t�0�1HD�Q�w��1�JN�;*���Y�<=ɻ/�n�Zv��{r��Ur.�%ߌl��&秭r��]�����7�����Nƞ{feUe-d�,Rܩ���D5��V��{�16`c�c ���6�M���0�L�[ݒ(Q�"Y$k�ܷ��#2����nf0�T���.�t��/�{w=��|������=�ګ���U�b��ŀ�#bU=r\�4�/ttGF�!}��w��sz����l%�M܆1��e"A��t�W٤Q��	����|)m��EE�y\�ZKv������0�� �<�0��b�Q\/�b����:
��eP޸��$k$O��$]�#�G	�l�L��}��E�E:��#r��;��Ah�������q��ԫ�q�$�����u��U؎�C���!��)��!1� 1|�!~�I>��{��czǣ��Cn =|�>�$�)ܧ
�KB*�����ьlF>ǈD�SvQGE��~c���z�8��D$'qb��F�g��_�>��7򜰌�x-�D4��N4x�G]�tǳ>/��ܴj��C�4����i8i�R��&�S�7�"M�F�5P�h�Ӕ��_�4��A#"}�0�Ñ�x�����I�>|`�N�zղ�f��W�e/��kv���6)�H�E�p�f�q׽��翩2� a	I�I�9J)]��������c($z�dG�H\Y��:�����AǦǊo��@�tgl�����^��_yɆ�/�׵)�e�O�����,u��	�p:��|I�I�6�gq��:��眍�N�
������Q~��3zb�C��GG�����<������<��j�OW��u�cW] ������Iy�?��
Y�rwr�'�DY\�I�R^@2�'�"{��tT����,Q>��l�ը���I����%G�c�u��p�[�i�5�y�����q��$=R�(3��~�0�B��l�ǑΙ���^d��x>��J��$��j�5������@����CĉT���L��<��]����}��)���i���ʙ3�#m�k�$mq��*�=�rPW�o4�pdƯ�ҭu|{q����ݻw�:��74je�7RFcJcd��5^QT)��;~�3�Q~ʓz_R�����a�����n��Fk �����o�o���/�������]y���x�C5�Ȫ����at�T�G�̣���P$�J,� �S��1�K�E�DH��2�#��8���=:�t�Yr� {T�W��ގ�����_؝�a+Su��M[����|�{�_��O= �ꗜ��
�<y&�zmAd�3�8L!�B&D���BS�R\��?&a�/ʁ\��q�*p݂hD=\B��y��"]8r�i6T�/�]Q"�K�|N��cΡ�S��h`c�'o�K>H�?��=��n,_k��^���:�t��3����.��E��Y!�A&u ��q�
{�c�SZ�v�,9�-����L��#�&Ag�g�:����9���]��}Q�@1^���O�gӍ�u=���P�P�3H�{����8�k�7y!�ѝcO[�]:���Ë{ "
!��z m
d��!T��l�|���:���I�s��9؃�]�SH:S`�yB:&��-+�f��#��e��������Q��������0㎈O�鍎�&��gǯP5�Ey�`h㜆�H�;!�1�_j`SÇCaR6�(�x��pg�����۷�:;m_}�U{�+�X�܊5�n�_�4�4�����q���Yx}8G%�M5�������3��)�O���(踝wG+Y�F�Ɲ�JpBA�WW��l������/���Y{�;ߴ���m[�v��""��b�/�Fp��3Ґ�z�S���8��ڻ-��=��S	��q��u���r�q��F\�G*���/�0/Ti����D�>��(�l���g��l>���)�nțKD�*��(�w����A��D��G�ӛg�c��q�-�	��#�Ħ)M:�ʉ*<��#����Ӡ�$gJK`�8!l�.�E����'�$[x^}ȕ��߿��{4r[��^W���5�ٻM��}܏�#6���@�a�c�ɧ�i'���0�)����t��5���I�$c:���U_�ǧ(T葟�eEy�~��D&��xR���ld���@m�7/���5��1[Z^�em�^��������'�3ў
G�~�Gc���QM&��NX�q����w���\3��煼8��^z���t�Z��V�ƌ���i�Su���(�2������y%K�M8i`I�H4�����U����cH����HU���vapG����Y��D8+5+��g_z֞��W�|aņ"�=�Vy��H�W�Q9�K�XA���Q�dDf�gؠ�w�B��>���a�&�k�Y)���@"�/zA�&����Bl����*vQ�ꆈa�!��J�~����� ;�*�������[ԁ��c��"��OH�|R^±�{�v\ZQާ ��Q��r�☼QO���#us���@8yOd�4�f������_�%�%��#J���7�����~�8�~*-V��RE�(�p-�� W@��K�8�	��Kq����B�R����=,��+���ܿS��ۈ0�p?AV���[�$��.�YX�w��|؊/�ӓ�!�K�]l)��>�v�'l��ہ<������yj�hl��ݵ����~a!V�fAP��Ј�k�bn�E�u�2�R��2��~%BhtqJ���n�m��/m�ᬨ�������l��e�.֨,��2��WhgF�85�^�WCî�W�ֹ/�J�=M8�h�C���_Q�����@[�.�0'hғ9gN��FPFaϧZ���ϧ�l0h[�3�õ-t{6sn�/_��e�j��]gr�+]8DOmG
�=��
C�*Wu�t!Ky� ����;C��!B�'G�D',p:���A��I�ΏÞ�z�:;	���{�T��n�t}\+�V桸�[1�; �a��zx`!'��8���#�:�(���'rG1�,E�p�\[�1��Ӂ�_T��Aa�a�v�pꎲ�A:�,�}�쿊$K�	'�_;Ėd�8��9�+q��⺜F����
ϫ�~Os�ci���k�׏݃��#䄉��3d�C
�(~@�.����P�t���y�S�4�J�x:�s�B����
YB0i���\����u\�H������ҥr�ǽ|��ۃL�2>����6�}юFӻ�uJ����X[[��?�؏gf�j�
g���,z>�5c�,�7�0�IQA�"�įX8����N��_�
�B�x�*�RM}�|/Eu[�.��nE��c�F��J$�tQa4�j��#���G�u�p|��G��r�~��Hr�Bw���a�Ǧ����~����S�8jz���c���b�T��Ϋ1U�٣�5D�x��aI2T��J���<*�I�6���	��R��%� �C�-ȉ_��%��~����@nő�D�(���O�	��q�% �2I��$}��^�QB�|)EH�!3)�:	F��IOQ�k"y�*���$�����I�c��8DV�CvB� qmC�DFR� `N�.��O��j���7H@
R/N�A�H�p�e*^Zyܧ�2�ǞL�����I^��F*��^y��㸦����CrT��
Y����_�S��d��i�N��3�	�"��GU~_7Pq��qm��M%Q_��ޛFC�|o��N�K�Ơ�jee�ΜY������z��G�'t;)/*uA�����|'�3~��IX��O��p @͎�i���|x��޳��-�7���w�h�u)����bœb�ȹC5����#�@#D��O��T��!5rx*�I���7e�w)�*",���!]�'9pܱj|�3;�Y��1y姁'_�y��*(���_�C������pv�,��B��Nӝ|C�	��#�5z� `d�Ɂ�^}���L6���7�r�⯰�G����ϑ��'8�e��P9)�/�����$�?E�aN2U��)ٰvI:s�8w���*����H����ޔ�^�I�=G:v���ڜX�=�:B���!;v��S�^<�K�ʢW�'�{MJ�r\!�[�x�IOC"��>�&^I�+ǉ���aG̸����M�!VY�+�p�H�|�T��)�"z�H{��<]�����Dc�$��=ű�D>�O��q,����S|_x����2|���V���;\���n���ں-./�ًlZ���vT�@�B��ߨ��ŅE��Y{$FG��T?a�C��-���<l��1�	����/���/������WqRv�k���4��2~��IX��o߲��m���:���z�Pј���pz?���xxC�d���O�䆞~�dI�#��Qv��!G5����Y����O�{z�8�@] yS<q8C�T7q�����y����9H士G�����O��(P�Ce@te��s�d;��D:�((9��°	������L҇��������K�A¢�$t��a��5�� Ɉ�/�����4��m�0��[J�=���9<C*� q�)�G��;s=�W���T��N�J�4>'�ʺ��PRޟ���d#�
;*�)�є�tb���	�čs�GE����,�/���q=�v�]a��Bw��/�FH�x����dTy��*&�)�Դ���C]v�c��N�G�捛6���Fk��޵n�Pd�m=���t�.��]|�%��^�֨d�A��Jy�I����^�[�F�>�I����⸎\ߣ�B��6~D�
�3g�����s�w�L"����ݦ�G}�=������wPF� ��^�k���hW��~7ӱʹ>8t���ޣ±��N��Y���׺硱U,$�8�	�"ՠ�C1)���w"�P'OEE�y���$ȃsK#
$$|�ىa$�q������nI�I�39��֑B&N8����1d�_� �["��!��	5H(�a� T�K����!:��QN菰��q��J�z Y��d�@()=zEV?��,/㤜@�8��.� Y؏�aO�I�Q��}���S8e�دe�,�≾�	$�\o���ѱ^��p���/���JV�qU�Ш/B"�2�˃"a��$u�k��T��t/ҏ4Q�T�z��$Ƶ�B��P&C���xK\;tKi�]*P��4�/l>79�˖�*�y����3�?bT�@�;O��D�F�'!�SՒͫ��?{�^�7���nݳ��v|�|T:���Zgn�ο����h+O=c������R��,)�еĜG	��J�mCO5Z�m ���C�I{2����wn�����i���4��I�#3���a@P����5 ��M2�c!Wo�ժ2׋�xqn8o����ڢ��$��o:�=?��n8�p��C�D^@^��c>
&�z���^G�˃�IEC\V �H�*N�2�h�#]*�&2�M�Cx��g#��H�R=HaI?O�sO�c6Ȇ��QN�Mi�)!lC8ez#�i9V���瓈�R�E~A�F ����86tI�n�C|�O�Ov�-��Cz'p�O9\��Z�%�I���2��aO���Bޑ�	�8����Xٯ+��"?*�F�"��&(���ؗנ��a{��_}B��5�C��p��+<���$N߫��~�v{>t���-�"��=�Nɣ���ʣ �	��wx����i������]۾����m��V�'�a�e�ۛ�Z��0�[Z���맽s"�n�F��K��XF�'	�7qߒ1��5��������ഭ&��&�l\#�_�7���e|!���O�#�1VV���������]���wR���d%��dC��k�U��Ǌ��a
�V8!�)������q����E�u=J�M��HD����{�8 NYepN�;���p����!<B�M��p� ��-T����<:�(>
c�|�MiqE�$��#�8�����i��<{@�p��a�<����"iC���8jL6���zcs��-��� ���>P�����{ot�\����D���������1��_E�T��B�{�C8fh�'�Vi�{V�Z>�D��3*pl�!���Rݪ�cp	�G���N����*��D~m#;����{��[�D�(Cez��Uah�	w®��X'�Jϐ>�~�SU��9�g��}�z�l5�]���vӚ�kv��n�}�O	"��ٜʩ��z�U��ʊU��T�A�j:�T���K�ܒ��B� ݸ|��R1v`��_� L߯ԓ�9i&�ltb� �e����t���$,���ХF�����]�p��f�$�M�`��>rB8�o������gʖz7h�S��F{zgpnN|�06w\*�:�,�|�E+@�QOj�qv.P���Ty NIg���x�9�)�����J{?�Ϸ�	)?8N����C��㴑P��\�P�N��xM ''���+��M� �@�O�ؑ!�ǵ =2�� �Q�-�E|�O�Y�Ka.'g:IN�y#} ��&F�"�*�O�UE��{SE&b�L�B��/냡u�6���]�?X��֖�ڇV�hH�i)Se �P����r�lnO��^��D6��d%eA���w&Ż�cW�O6)M
�{=�D�A�-eÈJ���c���Քw�\��ۛ�����hi8��R������3��g������7o�>��j��}Y];=;����1��l��9��ϊ̉4���_1D���B���q]�X����ic f^��b7�l!s[ >ᴽR{�ʙL��򜰌/$h ��+6�����{(Y�bss�h<g=��s��1�S��`��,f��$���S��y#����:�z	'-�7�|pnj��2	8�TH=a'd��S�z/�^/�D��x���8I'@!�Ic��h:��4���xT��8l�C�iȍ _�I �����S� �8I��i�Dq�v��a7��	=�C� ���ѕ�d/���܆�q}|S�QF���Szl�SmA���u,��$�δEٞ��
��5	�� ���?��*<z�ƾ�0a bU�U�hз���D$�߻i7�s니��M��6�<7m6Ӱ+�?k���n��%��ZO$�;�"���$]���'���e�?�)l��FA�'��	�N�t�2o
"*��$��^Wʧ��i�%�Q>�=Ő��!��n�O�{6�������ڷ����x�ߕmk|e���܊��S��]�=�}�<x`���7�6+��as�ng��{�O��]x�e�辩����~ދ-��y�A��}'y�yO����ȝ={�IX�w[�p��6�Ǿ	~�䙼����ɴ��{�2��H΁�,5r�a1D��=a4�[[[Sz9
�BбuҤ�9N=\8)0YO�E�덱�� O�G��e�6��8�S>��Ԩ�U�����^�C	w9S�pR^�ץ����L���yr
���*l@q�q���Մ='���{b��ce
�ܾ�r�<*7�5	�!�	-z),�{������d3�sb���	#>�BƐ#���+R�����)��2R��T��ОwM2n�-U����Э��K���~t����=|�m��w���m�枍�v�����������!�i���e���{E�DI���a.'��{�t隸܅'�c��q�u`�$J��y��.�f9����ڌ�>\C��tg(�tز_�����?���+5�6����TL_��T���l�-��9�Y]��k���3��zw�l,"6����ίڙ+��ܹ���%k�qU����&���sT�n��9w��|f��"���)H�I�J�=�v����{4}�22~2	��{�h�Q��0�`.^�sj��ݻW4� &��U���1����A��������Y�Ԏ��� �jq�DcZ4���|�!�<�#{���/�H��X�9�/��𫛺+�|6�^�a/d�B��"��ɺCGʔsp��`��.�2�zR/��y�������pd�m�\����P�.�@�p��H8�E�
��.")N! Ed�l�����؎=��9�'B�;ɅLD'���l���"�D�[SM���rѓ�H�Z�aJ/]��.*n�Z���C����`k�z��6u��}h������E�mkm���Vg���:=c}�/l@�q��{G�"�m���d��7���.�G����&������+W�a?���h`���*����ܱw�ßٽ�߶�(�P^X\���y��^��%f�뾱���43�4"d����C��f5}�Y�Ni��HDoqe�I_���Gr�����{�Uy�՗b��E���Ť=	�����$�XK[F�_�L�2�~�px����rrQd�u����<ON�(���|8���uBR����v����_�8���<��=�8A��4�!�yx�~�G5�rp|N�F�h��%�z��|��Sv�9������X�eFO�r8Oy��e�H�i .��,����s���8�e�8v�5b�U({�!i�y�",�&��s�RI)+�zɮ��ݶqL�4��ޓ*�e�F8�<�p\~�@����V����G�+��7l�M�X�^�?Yx�>mK",q�i��ֺH���!���
�i�ձ)ݷs"<Iɏ'������:v@�I��+!��4�Z��9�N��=i|+��J˽��=�0�Xw�{~s�vo�o��=b�N�F"ፙ�[Z���y��3e���|��v�ǯۂ��̺=���66��<�:��0%��\�`._�P�*b�����|N�t��$5=|�Ϟ�E��}@�H6D�D�>�9�_���i|ZXF�$,��h�i���~A�^��?R����v���s�h,!d��Ӟ����d�H�d* ���x#�[��"� ~+m	���#�$2�M�,��zE8�0G*9@��3a8�D$�:\>�S��F��8' �tA��+lH鎏�CP/�̲#���_�C�"�¢l�4�.C�,�I�4�����C��<���A���ғ��$����F���Z;)��(�b�i#^�xi)�<v�u����1�w��ׂs�I;�������l$�sŘ��^��N�"+k�}���gO���<3՚���v����ڲ�q�)�/�@���u�$�m!9;�l��Mq��$�7yy9~���cQ@"k��-+�� �%�l���ت���������oݵ��)��X���{=������|���ήm��[�-k߾cK�n�R�������XywLLV���KS�KW�����R��65+��I.��^�)_o���k4b�(ךk�z����,���-O�Mn��L�2��Hm���+��n����N�1� ��߳n�kU5�,�ʊ�^�CZ����j�U��k>4�D��Τ6�j����!92@c�y��p`q�z��C����Q"iBw#� ����"�$.y�q�-ͭ��D"Ґ
�^��Kr$���"m���R=qi"6�����{�$_L,W�"'��U�I�޿H�s� �^<�*/���I{�CI�����<�΃4�\��'Q"�|�xC����
�@"�k���8�1U����c3��/Sq�m�P�d�V!��"d���H�ڹ�귾iׯ=i�[68h:y�'�'6�x�ƴ�/.XE�r*x��O�)l%�&{�@�+��}؈O�>҄^'�E>������(?C�<��DxH��>���o�{������6uص��HT�oՅy�Y]���%+I�-��[�C����6�}�Zwn[�ӳ�H蝷޴���������6��d�����e���������z�m��>a�z]��-$Ú�+�����p=c�[�0��^���i��N~Х-#�WA&a_Xxsv�MKm"m����0������[V��iJzD����3��^9~PeRMM:�x�*gBxr�^����+F����(%�x$��/�V>'�����Q:��-/���D<��Q�N�����C��sȔ������%��T�{9�'��L̥�^�p8U�-l��q�?��y�/i_R��"A����,�|��P��Vφ��Z6�:��ֺ�޳�޶�mJκ�cT�u&sWk��%H>�&Վ��G�(�͵�$�Ǧ�*+���;���.Ri&�<����S�J��a+tU�J";*>U@��2�ܴ{?�����Oli�nK�g�ʐ����nYi~�V��ኈCce�V�^�'�޶v����nG������~n��.^������aN׼$�ѳ���5�����ɬ�d����"��)_�@�ki��m�]���#˼�U2x�&�ɼ�?2|(q����zw�>%`��9{��C{�W�P	�Nvw��w���<��a˪��ݻu�Z�[v��ge�r_�d_�d�"�{��ٴ����6o}d��M;�|�f�q^m~i��}N�P��k�����*��8:L�&ٌ4|wا�)M����B&a_Hx�)��־�n9���)�����#拵�" 
���/ᢡ�2*����8��Qt��vS���\��K�(�TV#�BI<�$bewDj������(1�G��'�C�XOJ���,|���NV{ds'���{}��Yp���P���8q��鎄^!����i��m%�DJ��N)�P'Gԫ�";�^
c_N��e��?��߷��ߴ�w�8߻a��[wo׺�6�l�!VmhcX��(�Pf��^cgٱTb�6z�@8I�F��9�ӸGBg���X9���dk��B�qbn)*S�k�|)���ܑRr���ڲ;?�3[����}x�f$^�ܢU�àlU��U���W�vydu�9���=۝����u�=;���ٱ�Q��ƍ�M_<��V�:��Ju�ڠ�M���8�1�ז�w��:�^Wt�w2�q�q�!a�%l�=HN8=���ZDxq�X���:V�
�ٯ��[]�<�߷�;wm���X�V���s�ؗ_�٫�Y�Ekk5_?l~8���oY_�kZu1n(BV�H^��2�r��]��þ�����ݴrk��t^��""?��}Ϊ��U֏/n���j��Ŀg�����W�������ǽ�W����)2	����a���B�C�����;�iL�$]�?�Y��p]j|�O:+��8Շ��,Uz9Ū�{zQFr$�/��g�s5�v4P]��\�I��X���	��{Ψ76�B��%�{�ސH�©�zS �p�C?�L����2�S# }�Wcލ䁠@&�"͍5������/lp��M�4��߶���uֶ�����e�e��'�yo��``�$'�R˩А��^F�O�}�
)�'��)��臹�T`���i�|9mIQzI!�uy_f��e�ӋW�o�}�v��ߺ���ml�N��f�lvv�3Va�����m��M��6��3s6;�=�p�����`gǎt�U��^��l���)�X�D�W�E������C��>Q*���>t<��C�]ӆ�+��A�þ'�|XV�䤸��{�k�z]�њ��{���}��)�Y�̼�>q��]��t�j�yI���t��@<������>�\���ڥ���uo�CG�sZ�؁�V��X�<o�{}�-�g�z¾�O��jγ������S�I��
�\~I��1�;R���F���),#�o�L�2~�A�9�S�l�:d����닱O+d�8�h�9N���t!���A��6�6���6��-o����X��'a��4�Ho��(��R���Q�w��
㯐�N��8�t�l��� �(Cain��8���Y�x/'�1��!/%��Jijd������6�vв���E��6�w��n�����UI����ɱT�H�"�*�Z]��VȬ�D$iG��E��P�E|�瞈t����\�̢��}Q}�/��B���wز�7~n�>����U�[�M��Y��ԘnH��ɞ���ڻ�#kmmۨյy��F[?�y���~�I�yU��:;��>���ب��~U����X�!¢�<O+N��3Ѩp�
B����e=A�$!��O���/Ga؟��X��d����]��CS�{��0�S3�ml��9[XYr�<7Y���m��]ے�����t�Y��6���G;*��䓚�����vV�z�~��o���e���v8*�H?Dz��o.B���ˮ�	��O?��yFƯ��e�ƃ�4Q�������bL�����H��%=[8�('9"��x㆕�Á7�8O=B���C!���1�1�J7�|�U�{�y@�8O���j�rr����$����D�<���t�D/_����I���cBg�|��8� ΢T�yY�Ş06N� "aӳu;3;m
��1�w��w�P./z��Þ=l��5���Y�'=���wJJ�/{�Pm�/����%�[��	隞\WҠ�d�}�������JL�bLP&��"S��v:6:l[���;�m�:�����߷>+�?u��/��LJ��=���7l���m�����v���`ݚ���ڻ�Z��=��Z$�����/������Ƿ�5^%�wni�D�c¿d�WjV��e2$v�i�?�;F|7�>�|�}���&�،|�Ws�x
9Ae(R9z��M�g0��A�޹gG�V��~�km�j���@�l��k|l[o�g���X�B��zC[=ξ���V������)�O)u�[�{xdۥ��������_��}�J"w}]��t�Ԧ]ߊ�s�j%�LD�2�~I�اaǴ%$�dd�m�IX�oR�	h ӖE:N�
�ä}���ǀ�1��$��v�<@0���e�RC��q�)�/wB��x|�m%V�3.˙�������`>��a�|�.m.��!l���l��ER9�r�3牛��|��*��X����HO�y�'�	O��W�c��&.�|��,�;Q#��z0���<�[[���c����-r:I��f�5��>�U�Ė�r�̥���>�<*��PYT��\>6��Xa#��g@q&�T7z�p֝��A2��F/�_O��:&��Pd�I����v�����w��ԝ�Ї��.��-=y�U�i��wޱ��;6�;��V�J��>ܰ��Z"����u�Ca(2�]�Y��y׶Dh�=;�=V�Ul�̲ۗ�R��/�#HI.�L��|�w��K�^�irb�d�8�}y�{L���d��77�V����6���is���]}���"����[7l��]�m)���"��Vt]/�]���g�E~������Ѩf�#����}����mm�+�l�z{��G`�a�U���C�q_�M��B����C�Y=`��d��ŴM"���������!J��LާW�ƗaJ�	���~�F]�%�0�~L�>^�¯��뮯[��=k޺-��C3G�������1��1�z�cT��ϱԢg��G��9��8�/�:I����� mQ&��i���.�M����,JZW�Y�Q��l��'Q3"� ��Be)2��.UmnzƦ����`瞹n��M�D4����{`���z� ����.-[cq�{�T��d3��<&�ӳ���a"�vX�e渀�S:6�����v)tt$L��{*u���ŉ���Ît���ۿǆ:�i�)�kW_z��]��'��S��*���"\��]��D��m������n
��Ҋ)�^��|}���*��V�A�c�sv��V���R�f}ף����`<����5׍���1qi�� ���S�q��>rD�d؄�W��I�X��x9�����%�Hg]��eXU:t�m�nYg_�'e�UWyf��4�v����:�M+��߳�����_���i��U��˺gdk'��������0��4wy���r��N�q$�>����"����
�nH'� µ��d�O"O��ao��J ���jЃ��E�v�=���oZG��;��X��Gv���!۽��6֝��g�<q\}�_ c���EE을Qa�?�M����19@�	}So�Ň�JQ<���t�t%�X}���F�;'�Ely��ō�_	;��r��:3�y8A6���'��tU��sO?e+ן�3"&�]{�f�0�-k?���Ȏز-��ڬHZG���]��*��0+L�11?]�����$<�u�!Kd"�=���:��p�ز���@E����m۸y��{C��f�/���'���kWm�������;�/�7�1�F�𭖕��tx�ү�!�Gi��Y�/];]���@��ʳp���.�ѱ,�=ZG�J"7z�#�2�]�PE{���5���﹡��9�
r"�����V�9��wla�a�^׶�[o�� ��7Ƕ��-�>mc�H��Z�a�rߚ���{����ݎ]���������'�Y]�vE_?�j�J�2��	���<��7S��\�XBN�E�\O�K��m�32>?d��[��F63/��b,m�9���4� ��ي�Ͽ�F�}4X�����nӺ"�o߰��[yk��͖��d;��2bV	'?=U9�>�FN�eb⹻� #$�C��(�E ���|��dCN��F/��![8ϭ�1<��	g�^E������3	�cM���G��C�|����[N2��潧�!�١W�!}�d^���MW�רZ���(���0�9�S�	<V�n���˶r钍���'�(T��	����!h���#.�g�@�@�pN����+�Tr]�u�ݝ<D��m�d��HU�;67(�ܸ,MY�5�u6<+2r�#v��ܻkÝ};:l�
ٲ&R>;�5,S!�|�U]d��G�'��I�)_犫9���%�lk�sVў!L����s_��l�8pr�sz��{�{-�@`��E%8�rx��M�TB1ג�?�\3�Y����Qɺ�>�D"�߷�td�4�1P�MK�#��V��=�J�+��������e��d}�����^e��*GUJ�olq!��"N�2I����]��������<�IX�o=���-/�0$���W�U�#�ם࠘��0y��xí�%9�$hWW�/a�V�5��T������/���/M׭67�:��"����q�(j����?�T ���@Z��'$ټ�p��D����:�b&^��3ҧ=��/'��e?-Y�;{���G�������ذ�wG7-���g����Y��`k����OmwkӖ�.9�wg}M����v���u�Fҩ!�v��6����<(l��
q����I{�P��t���p�،�H�6�Fz�$}�C�aѓ��T,�NJ�\,ֻ��d�����1in�8K��{���ӽ�~t�n߱��C�:1���2e�=y՞|�ueÃ�f,��Z��KJC}P��x�[m�
�u_�".Jy��E_��hJ��*�`3��v�:��'@UB������#���a��ׁ^W�U��*=+�@[�_��zC��{%rz4���,N3��H���֖����;o/��?���+���h��%ce6l��,b\f""r���^�ҥr��| b苜�6�N��.	���2	��(0��:��y�c?����K�����>9n�'?ǲ �J�fD�fTF�i{����ٲa����V�wC$lj W�_���N۬��P�"|�ʡ�`;Ǥ̇U_�\�>rf�L\�G�J���Ȉ'D����x����$���
a��|��$ܜҵ�޷�_�k���ǖ�E2��H�G��UgglfQ�s`�����{v�o[��-Uk*C�6���{�6:ص*�?�͓�k+Kv��TC��`�ů�&;�a�) q��S-H'\������&�4�%xBi�gR����*��!���u�yZ=G�����Xt8Xs{�Z��[��[6�ڲ��5��iƑ�Dφv��e{�+_q����`Я����s�t�!#/�즈�M���U���X���0�Y	Z�
b_�Kז�������u!a�R[�������Gq�I��"@��t��gW���ܶ�¢=.�y��U�]]��+v��9[�����m����=,ٳ�}�����ؗ��?���s����G݁�cn@��T��cz��9Ӊ�'`�	���3�����_72	�Ș ·�w�hpL�d�	��Y�җyps�<o�ȉ�yU�6��`g.���g��V-Y�V��v˗c�[U�*���J?�mXi~��",������;��)��(�!\!s]�g�pL�<Ù����9�p�@/Έ^=t�I�^��;�ex.�p��PY0�99�死N*��XM�4���lT�Xe~N�r�fgk��۴�w?�͟��z��u��w��pݶ�����߆�(R��?��⼕�m,B�ps��y�-k�؜]9k��YL�J"r�3YQ2�/�=�2���z�8W΃XDD#zI��S�뜉��H�|�XĄk aI�ghm�V)j[E�%�k"V���z�������6�ڵ�ή���Ɗ�"}��q�]y�����H���<�0��a�ӷUٶ,�c������s��׿a�>aG"&<$��{vBJ�/m�'6	�t�#*�3l�g��	��ܣ������;�>���iC�ݮ��Y��h�ng�_��g0��C��ضuǥ���?�s���6�ē"�3��8�^,t[�~���*/W�j� ̅��qe���!t����|�22>Od��1��貟t��)�3Ɠ�����a�676��|$^�,"��!ӫ��R�-���Pmy���9.�;o��y�v����,���{�l(|zYI��H��,n�(�˾��rO酜8/z� T�t�_Ιyd�@Μ|i�:isrA	~���D�@��������H(�z\.W�u���ߺm�����\��em�f�hW^~��/^�������Ż���7���g��C_���w�mtx ��l��9V�i��՗fgm,��^KD����^8o5��H�,c��yO���t��HrB�9��>�=Q��y�W a'�6#�2lh-����<ٓ�{'�HE�h��ۜ�{���mS���*�i������<Iɰ�Ci��D���Ve ��p{Ϛ̗��3H���62�Mb�n����._��_��]���6�zVW@z��l�>�=�\3&���ck�C*����6�p����0{ �S�����e��w������JÄ}@1�#ŵ����`�v��v����轏l���w���V�_ڹ/�bG�Y}x���t�2�rz��E�w��O�g��ZG���M��T2C8[����yF��L�22Na���8m	4��1D�,����g?�����`�KglaiAdLN�ޠrͦEت3�6%Q?�b��3v��E��_��Î��(��\������-�^4�<q�y1t�%�;����p�ޓ���)�����t�;�pT�HΑ��.9_wh|R�v�� �r�&@�z�U�"Gn�g��u�)b!
P]��sO]��_��ͮ^���``�DX�Z�ƛ;V� L��i�����W�a�)�4��<���M_¡��ڑH���t��L�.���Dt�ݏu�,�]B��Nܱ�d�8�Sz��"�����@�G���KUq��՗m^���۶���E��&�s��q�xr�^����i�C�e�l��YK���@Ⱦ�DK:wu�\�`W��5{���ou�C��d�z�H�[TÃ�������!��c�^b����p��Y!K
��Ut�˵@HUṾ��(ǉ�������^ӥ��a�6����枽����?��{�[ߴ���R7��2������P�/��P�1D�lJ�P��8�6�a��xD�$,#�W�&9��b��{̇*�r��x/�|�'�ﶬSY�r�CM�K�6?��ޏ��m�no�4�<)֗۬�mfy�Xx�3dM����%s~� �ӓc�� �|�9IN=9>��������|_8!Sr�^>�E��G�)�s����`0�
S��mk�$��7���w(N3)2y���V_Y�����,5�y��u�;O��G'�l����b�dP��u�=몎K8�� ��^���Zq��=���z$NY!�Ő���Fh���IK'j!M<�D�i��	
2�-Mb��D���H�p{ܔ�%#�W�3}����f�g-�NuE��9�V],��gȱ&YTr��#û���HqՑ�c�0��^�hW������k�˗�@u�d�Z}�*�;'��+ի��t��3��*���X���ʨ�%z����}e7?�G�l�y�GBec�d'�t��=w~վ��ߵ�/�h���=A䞠.�b��o�t�}ؑ���w32�h�$,#�W��3b�a���W����N�*�59 �q����c��[�z�!�ѶY9�3��-)���۶���Vj�}����6��bKλ��t���h�c���F�KN��0��į��ip��@q<������t#��N�8IB�Yr��9���GCYdu�V����k��-��)�z��Cb8X��i������m�l��=�tdN��NP�3��y߇ꊵ��#��D.X'�1%[t�a�y���U�_�a1U�����h�;g�"�.�LpL��;>���m�?�+�c�[F��c�r%� 0��]^����m�^N��<Dh �>9u�T���v�l�k����t�y
"VUlOv��>Zz�Y;��p�IkK���0����6hF��Q��L��AP�������N/T��?t���H��9v~/�'n�^���SylD�7�:~��$��%��X>���Nï	ߟ=y�}�48Qf�[N�pdJ�_Td���7~j�!"l��D�!���y[:�l�"Z��={��v�����߰��؂�A�ٲ��=�趍�v�,�6��g�:?c����Y��y��S�֭�:���P�ɷ0TEo��ڧ'��ω�pb��A�	g��z�ċ��J86�r��|�W]�.����HSz�7iAz��M$��@�t��K	ҥ�* -��  -`��AJB�������m�:g��޳��<g��%'�U(����z{����BS�N� &`fBUd�m4���z�E#�Sg{wV�sl�L���fc�2�h}$Kkk�l$At_t�O)/v�pґ���y���Ak�*�r�ɶV�OBi9%��׮*^rce��0�-�i�S@�=�������5��.|[���a[)<L%S�?���t�w�l4�7ƒˀB�){�_��h=@���	'�T�ⳬ�m�'�T�=�b�^�ޝ������ҍ;i�K�%}�p,�i�߄u,l1�#oS�"�D}��t*X���8���_e��P7�h�G�
����e������H/D��]�%�������M���;e�����{QY�5���Y�����0��	[.wѾ�j�c�O��w3��I�d�^w����z9׳�����y:uF�]4z�ϝ�I�NK�N�s~�MpH�W���ϢH	Vc^�{7�p�Y��F5�#܎�j
�Ud�ɒ�!����*)x2�����4=����ԨA�X��O��߫��YVc4v�8z��f��RUL/�%�M �������{�&���E���P�ػ��� �۰���C�NpS���/��|ѨM���2�;_ȭ��V�t~X.��t��XR[��8į�VB���a{{�]Q�/��\W� ��Qt�z�|�P���T��14E�֓�W[�6o�_��g7�^4�JH�d��kX�o��xK��Z�ķ3j-��ul��Aȫ�+Y�<��dg<ú&"vRY1�g�r����=4��%v��l��ɵ��v��'�a/�5n�Z
�ڑ<��0*�P��z��e�+ ��-:;E��.��υ�g���8eD�������R���ic�Z#������`�����YYl]-���L�-D�S��\�۞2Dg�M?��2�Ё���e]�M���Z4Uz_��`�+ �"���Q�Xp������e��mݭ���(t~��W_PJRw�G�ߔ�]n�1��p�����˯���I��얒�"���N�$�[Lq�S�ն��9�� ��볮�G��&��:2Ԥ詤z����&��m�*�<J�U���i�otl����pQ"�$��,9(�G:�=x��: S2
?OD16r���+�^�,��l
��9��|�~$�Sڮg�nt�$%^���O�+�{�I�j98���_�^:�Y��.^�aU���YMpZ�̈́�ZY���n��-��k�z��a���F	��[c`�--D���N�����8H�u1���m����̨��f7�F�ɻ�Z�l1^�\��	ϔB�[߿�0�O͎u���3o�Փ�f8?l��b/�պ�*<�������9�ʓq���66iO�gX��_�BF����H7�1��<�����/�",�e���� ` ����h��dɨ�lw5z��B�k^ڃ�����o�yP9���{��e
Xj�a��H�F�,U����}N"�����>�t���k~(���\�3��w$:�6�R��>��d�+-\W��+x����o�-�E�/�����ik-�D���Σ��_�h�Ӑ��Jz
*�z�c>��\���Jj�	���F��o��W�d�
�ִ�A�.*D��ɮ�	�-6"�)��б�<�,G�3��Gč�6c��UT5�ͧ?e+@8��['��� ��rs�p{������cZ�s�3�T����E�~��4,p�|��,7�8I��~d�n��V��:b�\]8�H�m����,�y�(f��?������߀;����Q�	YL>��g#�@�>�N��5�F�9��,Q8q��ў+��(�_�g�<Wj��ObS��us�	���c���������nU�&��[��gTe�=�`|��z@�cy���fө/�[jYx����q���l�-2��Y�K���u}������#^ϻ�i<������G�D�JK���<�(� �M��=�u���/�!F�z�PVEj3��=��>�s�O}��[�^E�-��4+�P����9�7�Y������!�= ��4���R��L����ۀ;۸e�\�n�d����p-=_���CI�v��������,�������N���Ȧi��� Kl���b�f��WL��6nB]4�#;�dpurV6�#�;���[Z\�_��!�@F��G�b���0��2�P���S��3i�vy��sr/\��J��x�w��������Z���8&�����ܹ�$p�=[���w�İ�w��bt�������m��1����K��Ȩ�jiԼZ��=������s{��&.X�ˬD��p~*���!���e>���=���Ȇ����}Ow�n|l�_U ��Wj�
	q;{��X[PaT8�V���o�*�m^;{��2a�G��^��Se�Ĭ^���@k��J�����5i���1JOJcF��BŐll�`�t3���J�2Ga
JN�E+�� LP�ؒY���eԧ}��ֱ�O�d<qFa��v_U��G�8O���W�J������䖳��M������l�)J�������4�Nra!��L$��p$G�0��o���Q�����
Ϋ#sDj�%�&E}���|$3��m�������{qw]nj	)�.�*Hզ���N+F��hT�R�_,.�d�~�e.�Opn�Ar��af��^<v�7���e�5+�z�7�0�b�6��"�	Ѱ��h�!YV�J;�cX��n�fC�U�3�Xp��Υ�?^U�i>��݃�l�}�}f�eB�0�>�M=�%�_d?6�(������;�pg%[7��g�C��-,ݵ0�T�E���\�&���7xD=!b��1>�
s�V�C#�ж]S��U�x�Y����e��8촕���ȷ9CD+�����i�4s[8�Z�=�>o�ܫ���z�-1��W��m����G?�f�}��4�9����H��z mV����zI��Ufm�7�Dk��l�m+] ���7b��T�"L�J�H里���L"�T'�a��U�����X�r�X�f^���_G-�l#�8|���z)���-���;+ce�+H�8s�
��1`x�S��X��b�Y.��P��y[11E���[�Ջ9�	cX�x?�rK��#rC.EZC�8Z����Z�iYL��zC�����.Q䍕�F�e�}[��ew��L������@��-r<��Q�c���d^��F�y|�����2�'�2&��m��+�ϣ��.?�Oב��8w�ݝ#�Ϝ#�zR�������t����u�Ew&�n�w�D1]�����O��ނ�aOOy��ߛԝ/W� ����9R8p���r֢����	.:]s&2�8����v^z��a�4A�k�F�r쨘���������ꅊ�s� g�7��B�[B��v��:�g��~o��K��/Ni
=�˦��r[3_�=��B���*��9Z��d�G�����4ϥ���F�o?�R��}�s��|���ku-N�O�S!7>�i�;ʃ,��M��g��^Z=�q�i��������jx�����͕���Wc?�d����Y�=8�"���d1�����_ؒG�'��]#BT����r�xr��J���Y��:�Ǣ��/��e@#�7�1�#%p�Bm�`N��ؑߟE��8�%��m;�KS��w�:"�`�L����yj�0��o�ړ�X�X5�=�+��[[�������|!W2ד��V5��0щ��e�F���tK��tթ�5ծ��\�����m>e�Gs������w�\��X=B,%eK -
��#1w���8��rW�sE��Z�RK��7>ܘ�w��(GBj�n��t��şܦ]��K���z�<�
^enFwfȔ�ᡆfuvhP3�d���\��Ӊ4q1���1��s�[ox�C�����K�T�m�k���[��΂sF�6b*�ek.B�KqG,�2����O��)NH��\N��W�^�t�ڞ�8��VEߧ�MxÞ�u���N��u��<6�c'P5.4.���k ��z�v��gm����-k'#���]�(ȶ�L<��c��ɘ��2�V��A{�Ǟ`����Ek?O�#�����>#)PcI��CX�e'�7
T�+�F��oslm�-��ƣ�E����x�,��<m����}d�N?v�J}^�ۅUE�H�L����j#Jau܈+��-��S#cr#��l��9Sa�3�K{���O�2�̔�&����+�t%�����rMP<�Sߖ�A�G��V�RX��}7!}�/�ы(u/1|Z�+�0V�Q��B�:��e�YL3k�K_�Y���uF�sT�Ns�kLB��>K��-�X����~�I���h��R��/<&�i��\�O�&���Hy0�N8�������|@��ZV0�|-�l�ƭ��3�x��0�tm9�K�5�f���,vyhD�P��
b���k�h��]Ko�^/[4��F��V���4��S��Ta����A���,���8UJ1�p�eW��uǇ�6,Mf�5z C���3���
_��@m�#��2y��,ֹ�gP��0_��|c?|0���8kZɮH����<�נ��U�c��R�f��%��/��9�e��*���Y�w�0H:����h����%���	[��8�|(I`d���D?��=�'7 Q��?�� �R�ug��:"N� yNz78�;콈,�`g>G�SB^��޽{{�lR�K�L�R_Y�`�`+;��1�:�$�B����(]?�V�W�E�8�<�&�l(�7�Û�]Zə3���uuN;�|�j�����(��c]��O -X5�)��!P����]׎0����E��6j��~uI�3�g~t%#���׌�֗�	�ƾ��ϑ��լ���!�:�����0*���=޵�9�x�rI��F�n �	h����0;��S�{�(�'�UL��l��$��i]�ڀ*���������R�%�0�|�5�|�d����^�_{��6�)����~�[�f�7�����(W.�;Ԓ�2���@'ҨA^BB+g�+�ٙ*�PpOd�yT.�?�4E4�B���&��jV ���s�O%�Rn��v^���q7\�o�����L������_	�kE�b�J>����L��Z�%�&(Sώ\�]|:K��|��M=�ߢ����391���=ŷe޾�� J7�)h6���K�g�-\�����e�.D���N竆L��M*ߙ;�z$�0M���{mg%��������\�Nә��v�\���P��:{e�*M��E����{�{1D���6���_��D]�c��
�>	[�}�F�"K���r엮ɑϠ��6�ɦ��,?*�l�7z�ֵ���g���J&�+�%�~�Asm���D�d�ὃ?�~7�?�2~��:`��Z���I܊��t ��r.x�J�mP7�~�[\���N�Ւǵ��ȥ������FP�t9h�0N���jo��b�)֊�쬀�Tt���'�^�A�FJ�ڰ�t0�о_DZ�Q�F1R����]���
ͫIW��,Bu�W%��I{�������n'�Q\�=�p���0�}ni�F����\Ӿ9�4���Rm0nHK��H����Ԟ��Y��	]1������i��Lf�#e�"�A��Z߆���� �Y�5���X4���֫>�/���I�`����>-���.�>��Eo���O�m��S���T�p�i���J!�g�V=C��$�Z�vg�5!'{3��� �m�]�:�R��doYj�I�T�ǯ
߃�-$�3�~�$�[�C�j����:��eO����X�8��_
����C�����t��-�df�O]rPyЃ����7���ru�^`Նѡ�S���u��V���&��u�ά�z�����M ;�X�o�tK���|���X8�L@z�=����@P=%g��B|����+S*`{�wĹ`cv"_�-�O�M�9��M��I�0]�%w�����,��(�muc+�64~�n�����7Y��g���/:�JS�z�\���:lG���7Ɵ�^���_C�P��Ӥ�RK�U�X+���Ù��|��1�@B�|�����3���,�� ��&j����c#~�����:����/��\���q�&������)���9��_~���m	���1�3��*4lp+׬��܃
Y��Ʒħ?��z�>��f3������;�ʤ0)��pΗ_�Y��DS6��Mfz1�k?��%��b`��>^/v���˖�.���#�
�F���������&�-�[�(�$�Y�ˍ��_�\�q���� �.}��g�	���B������4����)w�����>p���đ��1���e[�8�Nk+�3�{�d��i綫�D�T&s5���G�Fœ�XTF�`$qRz�ܝ�+�I���9��|S��NVC~���F��jӀ��@vO݄��VD|,�������Źm���~�:T�Q����3�>a~
E6;DǠ���9�"Vxdh�f�B�"=x]��;Ȼn�u=������ *^N�}�B䘧[��]��2;E5qZz�6��'g�O�����Sa���f�=���f%��ov����IѴ�3��?�z �ݢ�� �����os�w`��<�wc��{��	�;�4�m����&ɰM�
!�2�VвK�uYZ^��O����)�R�o�M,p�����b[���?
��В��y�*�i��<u~�>B���뢞�la�ߝ��И����lf*����˕���SҎ齙of[� �Xe ����IX�-�Q���lWCi�v�!uc�|w`
+~&X�q=es<�������R���6���)���Wex�H����#��O��6�����z��ǥ~P�����f�wZ�0��t��	�u���-\U�e/�0�Վw�M:�kOj��n;Y�f�Sk7��n�\��V����9g�|?I��E:;8\z���*/�G�g]&�u����_1>R�L��o�����'U�H�8?�jE�EeDͦ$zzt�)�nH���O�=7�rV~9��d�/������m�jݟ���\�4wo5��EB��d$��H�eq�4Ȋ����֬X��H��qq��O��R��*�̱���9 ������9���:`@�F�?:4jl�Uk�8�Ű�EVL�׎#��8�]W��1�Ҳ����YџY��"���Od�ְ�;�M�+n1���_0.�����[ۦV��xfc���Ň~� =��1��5���"n�ԟ&)?�ܿ��?r*��Y��U8�AG�><֔��|[j���t�p>&��:��qܬ 3;wTߴ#��bc&�
5)(-��z(���)*}3\.�SØĜ7���U4F(pP�<�
�C��j���rM(�,� r�0�1�?{��d39��VL
Z�7��6z�W��M,�ճF�Ɣ��f�u_-bM�<��8��O��[��� ���W��e���ɨ����}47|�|Y}�/���w_���;�*�-�G����%�ڟ�����?H��T0��9)ŝw\55��X��yg�W��@��W��%��V���y���|u���ai�I��s�H4մ�6_9F"Y���#r��FJ:RC���=NJ	�t(��o�Qf�f�.��Jӱ	<V�I��41�z-/���Z�JN��h5�h��`Q�~�Mg��� �0�����2������]�*/_���-hd��t]�F�`h�6�y�K��*s[�z�[q������k%�~G��Xr�:�V��fۛ|�/	�|pϫrx��L�£�l	�M���;gO��7�ze+����(�8访���'��f��r���y�+!R����/i6�3�v,y��9����e�b0	@a��,6G�G_?�� +ys�$��In
~�- �9S�|����z��3�jl+�w\�z�]�k�.�'Νn����
FV�?Dy�����|������(��T@_+����3� q(��7Ru� 2S	ܱ����I��KK�X��?&ͤ'ߩ���r��v��7kr�.!i�䝁��@���vW�t�`���7���1Td�$�9�Tf�ڏ�{�dX�U_l��I-���2P3�ϲ��� $v*q���r�n�%e);$0w@S���9Mc�I�/вʂZ_23���:��?�5>��jL�L/^nL �����b�PiR�XkQ�:�|�f+I��%��'�l~In6������R���ێQT899!_~a��df��� U��ƿ �$�}LI4�������[=[h�sI��m5h���-t8�`���p%0��y�]^�X9�v�p޿�I�]����ݛ�%�p5t��8���P��#�B!��@�  (��}�Ɛ���Wkb'*�����`�9TSO��r��+�w�8�6�ߒ~��O�Р*�te�c���6`��j�Ĉ|�"���6UY���'�Q\
t�t��3�
Viưth���SN�������-2[�{�?�?��$+qO�#�X0Sfd�����;S˹�Or�A�kQ~G��l	Ӆ��0%�ؙ�#��_��혠�E\��5�ڿ��D��a��u�xf��l$��;#IK�~�K\#�R�)�}ZV&���yǹ��vzL�YoX$�D��*-�'� Y�GR�,�'=
���k[�"..�������D\$xL�y׫@�����:E�P8@;%;?W�v�;��X�T�%#3�8��e�6������C���/�M�����T.��⸕�nT6�D��25�T��[�����_M�J�U���@թi�#[��>��y����r�g�i���9Б�U�z}*�	���ɱ}_e�ɵx�~'�ρ�\΃q7�/2<�gez�� ���+�B�;�E�yKϸnm��(���	�R�֡��d(���b�+�<\��k@k�U?{�yJ`�;^h��#������B�A��.@l�Κ��M�e���k�u���G��KV+�O�>e������$1v���Ǜ��P��mG���d�ݙLFN^�
Ǭ6�r*��85Y�2������sJ���N��|�s��E��\�C�q����x�(�X�*���ۥ��>��i7�����x���)��B�g�ROR���O���yw�"�6f�~�PMZI�ٵ�㖿r�=S��/�vIJ<���O��d)�!��-��I�W]��U�T��}Pv�ԥˋ�h}�ؑͨQ�0��(���i�Ӂ���|�3G�T(�t��7�~��-�tW�I\"2�'�$�VHB7��6|��y&2�6:���G4t�f1_��	�וT}YMuN#�$G���E���*ׄR���{���]�م�η�d�Ȗcf�t�^=s�OO<s���Ļ�T�N[B�9n���k��E���'��lI�qю1)����є�;:��O�<�B�r�!Mߦ�h����k]8W��*��_�m����ɟ
9�T���t��@�-���=����w�?���^���MX�ƇX�qLZ�1�7����\�h��� PK   2acX�#�(~ I� /   images/e51fe3aa-205e-4659-a3a1-ad304791dd1d.png仅W�Q��=�!�C��tI)��t�4���H���J�t�tIJ��Cw���>�z�ᛵ\�f�k���y����	S�$��N�����TA _�*2�X�����(������BqO7x��UZ�U�����������拽������g��#2�$/�^�q���~�(~<�}�̨_�286
�=�<jD@ �G��a�nm���&lz��p~�r�а,��b�I��MY!N�HGO�k�/Ɯ���c�ܪ����E����)��U<�cO�v��η<zyt$ǞUr��zĽ
�!���D���h�r�0��jc������`Bw��d{���V~i�;<�٬R]E�Y���z���kWA��}l���3���gӏ�x����\����	�$	m�u)�Hy����@o>����t"�o'�������^1k�!��g�l�BH"\b߽�~�����1��O4х�bs���_�ч̜�Xc�2���kN#�Q=��
�#�[�e�Gl��V���"�#�Ü����fɬόzP3��hyz)�*YAPW/��	�V]I����')G6��������\ys+)��������R��F�|>�kb����p��pdG�E3���g�}���|k>{C�����8a��-.����06�<�t�y[謤���<I��#8	1L��C�~���@
�Fʩm3�9�oa�Vi��2F+J���K]����ԟ�K�a]je��Պ��}+O?M�C�P/Z/��o�fs'gDDmE��h&�1�^ۗv<��Ԟ��)�F��3�}���A�gP��w��`�y�]5;;/�)��l�(֌KKϩ�I� ����c^�{��&���ar�;:��nż5�#��ݠ�������a��3�v�0�s�� �\�'��Z��&�_EE@ַ��j+^/���_E�9��R����]�O=Rf�u�2­5��r�J����-y�&e��=��&��c`�G/��QZӌ��Ablz�k�7gU_2����@G�\�ل���߁�@�o�^N�y5w]�����l�~�M���X�:s�O*��qǁ�/m�3:P�X;�xI 2��r7���*i
~�W˲����͹�N5����<�Փ/W{U�����>�kv�$��IwU�.�)��M��6�c{���mR���H�����c���ʒl���&�}��<*ޑB;��ϑ���>g�.T�|�"���%��H�
ӦD�� zY���}���a���H<QZ@Ũȴ�w!/���?s)j�͒oa]x��oFh,������1af|~��K&�Dz�=Jߜ/N�m�ס�c��R�+��g/e�|�Vhck���y�f_�� �X�Z��酳	�����a���z��0;%0��ԡ�mXbp��r�8�?��u8�gvܑ0	��6����a��ԻGO%s��0��sv� .��@s��Z��=����;R�?� �=I�v�V�0|�褣��I��k��Q�nm)>sV�N��u��r5��Z�J�����Mk�p��I%#��F\�o�(��4P�1FO�3����׊T�@w4�9�VW�U?8lX���3�ί��-m�C��Zb�Ԯ1�k�0w�_m ��nq�%����$F�LO��m1�"�~4����:M��_N�׌v�>��_�	��7�z��N3-���Ъ �mAHɏ%uhw�	����LF[�,:;���	�����chbe;%Y��J$���0����G���Zi�Ȟ�m��_��N��3�V�1��xN_�ʋ��:p���=���`�&�3f�8ۢaN�U��e�s����;�8h��&~P���W��_%v��,��%S��b��X��࣯��]����������u�
�P>R�Bp��)�]�	���O���tQ����>�W948����b��R�<tL+�88�WFJv=��A؇ռ����]9ޘ�%H��P��	:}�0�~�n��5])}�%0Nļ�e�qC���.i���M�[�xqq��\}'f����V�wd�O_g�^�"/�>��� ���Z�flȿ��(�d�e��k�7��캆PR,9���\F�x(
˟�����8'��}�y��%��e�W����l�H("
,��'�MJ~[_�����"�"���Г?\�.�5H;J'BP�e�
}G�
ՠ�D�˽���%bآ�"�d�����8?�p������'����p������G�󇻰�0��9��1R�����`)������ �2[�J�6��k�~�g��իD��#���I��S��oHm���In�[!>��[1�p_;��>XBC�x���if��nrԺ*n.&$��F2H����،���a�Ǆ:j���?H��裡�e�w��X'�U��@vN�	vG�,s*eR��c��R����f���]R��C��X
<86M�1�'�=v}dz�b����Z<~�Ƶ��Jz#���+r�c�><�$�$f�w/���B�O����iԚj}2�.6��z��I���X�$^��W4�z�yb�~1�C�Nu|q�2��bBh�v�>��h�a�M�Ʊ_W#��fc���)�������'9��q��v�8L�d7�7:ƕ�d�S޴���Jw��\�����X�����7K�H�0T�����ታ���`<���H����蕓F��4)=�/�_�}g������f;���f��>)�:�Ü����Uv���<|�/��Y�L}+��ԛ�ѦV��Xϸ�8D�SZMO���(/W�[��췅W�F=�;�
`=�]k^aw�&���|�Pƕ)������L�Y�Ğ�xj���<��_�*���$���"B��b�Q�W��	���>�u�3��	�ث�P0!������K�4��[�L.a~|C�Q㙞�2��[�w��T�wCV����EMW?^%��<��5�sU���ߩx��Ʀ��H(�O����R�;k'�_&�>y�݄�Z�{~`��"4@����Mz��ۿ>���1=X��n�����I���*!��]6�u$t�1�oM�${���w����cR��{��#p._�ɋΓ���k�ӱq�E��=[s.�� \ܕ]�I��8������<�iz�������ճ��)<Z�:�Eu@��6��51���K|;�2v9|�x9������>h�l�Aԗ�?����y�t,t���tN5�Nk9�l����+�����0�'��p��$V�u�Rm)}�؂�0C���b�;Tz9��5�EQ�6�+�y�~�����V�"����o�q��5��|��"���>w�j݉PZ��S�FP�??��Y��T����aJ����:#�Θ=˓(��-v4����Y�oBWQ\�"?��5������7O��PP���t�,�ݏJ(�Wẁ������n}xɹ�g�_��=2�����E`˃����H��n�!4g~n�����Sɍ3�%d�"��EpӒ��:��Q���Q\1=��h��+���nM`V��g^h�4�i�&z}���)epzl�7mS�<���^�vG*-�t"�.k܇0������ٮWW��B@�����|��B~�-s�*�<o���E���f�^���xi��F��s��M ���òB�߯��4�}p5�=H蒑�J
Æ�ѼB�^���{1�%���8Ʉd�&�K^��g��1X{���p:q�b�(����<��N,���Q�t�ڔ;��I�'0cbMG�Y�¢�Y��C�U�%��BKȴ8�6�W�� S�$���{�/M?�1��˴U�v�׍��O��������߆�&P�6<�M���և�g�Ϻ� G6��%$yᘤ�C�;�^(��N��Wv�vZr���'�GāHH��L3�[�VT�W��D@2�	�h�˓�pΌ�6~�����XB������@�k�="��v��;��h�\4�:��ƫ��U����X4�0}��C}x��G�����9Ǿ���O-$��xɑ��H�?L�z�� A,�[;]S�N5|윱��);���@��ھ�6UG���X���
��fb����6l���߫AB�C��H�QZ��l�Ccε荹bؤ�K���e�8�2����9�O)��5��Q��|4+ytE"�O�:3�1ٚ��5�HۊyI��к��h�h&�̀'5�x ��1�f֘ܖ�Ia�~��f��7t��V��q��|�eU����k�،��*�[�}���ݛds���5Gn�q��t�.c�h��W�.�,v�Za/�"hv(��໐�2���be�"Q�l���V_x�=��Gv]Η?�@��28(l4�����j�>Ki�f���.�Z��C0opbcҾF�5�v����z尷>˪��a�Æ���<�W���3e	�ֈ�����{G��ct�b��ٔ����kQ6����pĝ��ia��T5���|���n:�}z~�wz����6�
`��>bqi 6Z%�X�V�<cOQ��/�NkϜ�ZZ�Aaic��&��1c���2�b�y٫���pX?��p�%%�/�E�z�D�]?�\��Q2�?Lg-W������-Y�۸U���E���Fu2
2Bd���:bͅ����eDVL�F��˸?��؃�r�e�lU��u��|o���q�̄ǹV�1O�������qB(��cT@ݮ��slhB�N� j�x4�쐈~��ZݷN;6���P�P
N���6�6���ػ��MY!��f�Y9GH��+E2,��ў���''�����~Yt�x0��w}�WN<�-�"$b��o��ҍ�j��&��V�|N��i:e5IM���J�����Oo��e��F� �p�׼(S[S+<ɗw��(���Ý%�~sn�K����ڔ�d�'ϽG0ñ�U�a�����+n�u����K�;:�b#4��MG^��`�?�����isӬц���w���]{�vz7��h���ټ%s�o�����٨8����GdE����c߻�=�N��.�>~b�UD�)�؎�.z�)ܛR�s��[���BX����m�["�G�h�=ҭh�s�o$��~�Q�B�٢�
'YLi{�@`W��	t-qk=��m�JR�٣�jB���/JQ�B���!����<�������55�k��O��͇�圣17^��|g��U-ote��Q��y����z'6�;�$k�L�"�ʘ�(���VJ��M2�6��)�;<kE)��p����cz�DaW� 3ǡ���,��#VH�5"E������H_���ޚQ�_A1����ǌ��4u��2yE���"�kM�V���N�ECn����@|�{}��Mo��B��LcN��P��Xp�W�7W��O{���/�4��U�nQZz��׈>����'
�w7�� ��|F �i�����o��s��q,�� �)e��p�]���y�5�犬�����u��֮X)������U>"d�$��Q8��T+� Yn]Z�u�c����er,���MZ @�9��~�d~����V��l5H�̲Ng�����U���a��y��cK9c
w/�B&(U�~،����	_����:�\F�6yUJlC�;>��w�����!K:E�D�(T���=C�k��T,U����Z�l�V�Ƅ)�5�԰�T�T5�M/?a� �z܆��Wx�~1���K�]f�H�nElO�5,���I9b��iu�5?t,q����r�{�؈��{fR0�ԑ��/��A�`��5�_�Uv�@��rP�I��}��N X���e�GVJ�p�#��fO~_�1ܟv�������������r
��Z�p�7;��������s�!nl�l�6�;.���04��'Ⱥ�^G'��qd����*]>�ډ�%f��6;攑��Ǐ��K���L� r�o�q�K4
��3I��#��I*k�2��$t���R�u�H_F=�H���f�heq�?����>K����;fzX�T&\���w��P���۴�eWg�ŃM�l,�_eSӿ�kZ�PGą̃A���z�;������S�P]<'+��7�5�ɲӧ%��PHf�0D�������l(�Ga_���v4�ZtN�hio)0����?������mfޞ�����"Y��o��7''�<J�X1޵�����AXE��?��鉷*��b��3Y}jw�Z_��2e;اК�^!^�"���A���W��a;�R΃�5¿�n�(��?���J�g�S�ו�`]�t�]6�B�/JNk�V���d����C?���*o"űZ�v`�.��f�%�=���u��S��r�6�T���� Gs��LNW�ig˞e��3�&��.�YWﭭ�r_�	�H�(�a_�eC�xPtJ�x뷭]	�rX����������1�Ct:?Fqdw:��\�d����*i'_x�\�"��6�-CJ�m�}��
䫃f2=��5���F���p�����n�Ѥ�J�\Kl���H>�|�ֺn��;�b?��!��c�3�C��h.Pc�c��Z'�Z�1�v� ̽�'�!h��C�����F�BVC'�=��y��f���b�b�) ����QB^j�eߝ]�>��{�?:�&ty��]u�EĞ!`6�"|�̑'��p*=�w0���k�+a3��E�d�T���z�U�|_��nU��\	ED�)�a��g����� �L�8'h?R�����e���0���`bz��s�|��Q���tx�=��EP'���x�ph�@��e[����4q���LN��!�
�z�6&�6Ǘ��t�mp�;nB����[�1�5s�R�5�-7�sl�P.�'n�m�rXl���7���=,/�
;�2`fW+Bn��u�m�RWB�;/G�H��5_Q2�i�[bD��bc(��B>������e2G{B~w�fOK��3\=ő��L8���xK�B�D?�&fwy�d�_�Ue�Hh�W�+N>�e��yZ�E d�d�<r��^ݠ�8��Y��u`�i���#l�P��mB�xp7We�L���@M�6�kUf���Z[MH�tA(�g���K�EG���=<�e�.N�!�nϙ!����L����I�X���c��uO3�)p��.�1$�ɰjc�T���B����+*4����q�Z�Z��m+Kr-�L�v7q����������Q��_o�����Ǐ1��u7]�uz��:���_*���+�A�c���s��F-���N� e�T�8����`�Ub��^�v�f�x���l�V>���t^�ݡ*5�Xd�m���g�ci|p��g��ⵡ�PG-Q�Γ�Bs"5���M$))�0zyw�;Ɨ}&���T����u�2{ŏ��(9��z�ޖ�eɚ�a��Ҫ�4L��QV�X#E��v�du�� p��r�⽠oT[8�z=%l%"{t}�2���+�j?-����w�޳��=_�{`�h¥�^hU����,����T��F
:����M��5���/��n:Ɨ/A����C�&�Y�p�(���b�R�o[�b�źwQP9�1�v�X������ә��`�E�������-����^#��I�#���N.�������R�w�`]�̅��ѓwDh"��-H+�
��s1��7mA.o��d'���𽌨UR�c<}~�kC�y��5��L����bh��߷�&ԅl/�DYtK�$JDg�ʦG��g��H�qH���8;.�T�\�3}.�H��������Y2_�LV�+���a	��ä0�Rf�0�+d����Ko�m}ױ��np�����DR+�v�j3�����Y����q�h��w+d��j��ҩ8�?#���p��+�c$��xѿ�<��6�Тڌ���6joy��֠���Z��z�x!�>I)^��HJ @|];�ͤ��[��[y�_{^�t,Oj��z(�W���J\�Pns��n�������4ZlV�Le�X�Q����a�Ox�KUy�p!�
��s&�����z�UM�&�jz�Z|�b�?�]���ι`���ú ;�a�g��]�#_�s]���yE�m(��2���.����[�/~�j�#a0���o��XO�Ix��.���v��[����?���0��Zí���g7��5�l(T��l�z��T���s�Ee�p|�Y�zxF�7#?��_[���bD��=�ѽvȍ/K��絡è���Hx���h�E�����t_�rk��R�9֡�I?1(�odo�^�^#:��ї��lC�Z�*��,U��}̾�C���Ս�6qsl��-��!�ۏ���t��$Y��9E��_�4�%<,]�#F�F����d�}����x(�?:S�݈Иʪ��
Q(�_(�,/����De���^�ԑ�-%Ev�0�P��ļ����a͈5͟��tG�b�hql�fb����������d�.��^�~Y��-��E��5a��ɝ�7*+v6��9k�����i�̦R��W����8��&j}�*��$;,Z�%IO����A5�W��b-15C3��(@$Pt��eĒ=Gō" ZI���YV�SB��=k�2@�]��Fǿ����ɍ14�;4������L���j��<b���|Yc�$�N�.K/m�EmBZ@�`'�p����>sc>������j=`[���D����d��~��Tt5������L���"��X�"p#�WV$q�}̆z��<��	�RB�n�U����'�q���X���;r�if d�ډ���P����#����%썺���TJW8���+�t�ڋA��L�!=��S�K9�5���4�E�M�O�J�y(�#�j���}#!h���������{,t͇�x؟�E�,�~�'z�C�W�:v��Դ�N2�F���э���<�ޙ���� i�S��-*�4z-�n������RW��2J�J���Ɯk@��N/�Qӏ=�l{ ��=�!�S*�-�Q�p�J�-����B�晏��q���ow/�k��P�t]ᅂ�;@qRl��s	�������⢝�%fcE�g_���;3�/.?���x��;>��k`��{������ϛ�M,_�@��c�����o��g�֬�*���6W��&+酔v�L�U��q�Q5�c٪�Yh�Ľ��+���0kV�˃�%V��ѷ�'���^�ھ���'�z)����#��b��ױ��`g!fتj�ŷ�Wvr#}$K~��U��MeN�,~S7�S�'���Gs�y�����:�/�To����$�m[�Æd�������J~��� _{f�#,�p*��$z�D6���-.��JϿȹ�+����BU�D���7�_r�3K�!�ͪۍ>����w��e2'^�۷�-�Uʅw�*�+'���葼���`B?D��Z�{i���y^(�cw/�^�Ghd�K��V�
�C;�Y�ʺ^���y��y~,�PH���e��OP�U=m�q�]��-�!�h#��+������X� �����'�=���I�F���"�k��Xt4d����5�'%m_�W�%f�ϙu�*���|�t|�]�{��o�t򏙉��Z���qk��dGri��k��͂o��ihg�h\3Ʈn6��S��q 	Z2!��¥-˼c{4��,������~�)�j?�j��eE�����C%�����z��X��K���mb���/Ճ��i������c�}v��݋�C������U�VD�"����?�~�3 �wɉ)��p�c�>��-���txl�E='[:$��bs#���J�;3LM�	��J��F�3)9�3H1Hh�H�M�!#rg�"�BX+��,���
��T�M��K&�QzY�E����|nhL�A1����#�@��*�3�"���9�����|EL��ҫ���	���G�8��l�^N;��R_�911I�Æ�kר�.���D����8�Q��㾁[�s�[e�jȯ�p9�>�-S�y��zű�-�7�}���b^۵�m������/̊C�a��*��n�U�R�<Q�gDK�A��E�� �Խ$\[��sjY�q���z(�:�;��	-�L���R�N-=-��	����(��!P�|�������s�\�W6*n�x��a�#q%�$}�2^:|�z��Q`釋�oaRZa��$݃�!w�c��[�����4Ծ��{GXB��],;P�;-������k�Ʀ���]lB�Q;C����ov�x��=���:�E�p�}����N[����˾��{{��Lfˇ�o��F��dzdۿ?֠��l������/H+Z	���iYa��:3�@'Gw΃��C"�B� H* ���t�OR�0Z�m�R����^t�
a[�!�؍j���ڻ%�D��Gl _��^'r�����c�_6�W8�_;��Xk�S� �K}�V�qg!,��=+�"}*���c���C89���eduz�_��z��E���CC֤��b/����y��9>=R�r�9�ܪ%�.�����=���o}�����
�d>2�L'z����� �'�������ǁ鹞��踜�&���b�T�plb�NĴ:�ё�K�<+a�(EUGf!z������r�Y����:2z��.�7 �B/K�:�]�5DkiסL����b��K���s������h����o
��e"J�O�:Ѱ����`-������T�I�s/�՘ypx�9�:�%`Nz����kN��G�qz�P�9af~�#gpؚ	��G$���(�O�vH��d#���T��CW ������5������(SkHP�dN�U��Z8����;�l�?���@����ª.��G��J�)�����m��߂�|9�]�f�*&�]r�JĴ�Ҷ�@��xPM����3��#o������9���$%d~�� k�DB]Jʾ�ۖw��au��۬f�qօ]��ߢr<�,@d�ʪ��ڔ,J�ʟ����{f냵�|��FH�?�D��y��ĆP*Y�9gZA�T��ׁ��r��B|��	�%|�8��iЋ�f�i��c�P:��.��;lP�Fi�TF�w����������đ�1Z�{��o�4�,L�-�\)���[�,I @A
̘�ޕ�R��'�_d�����[_�g$�plWc�rd�)���Ƒ3h;����]�5]��������.m��&�U�n�m'�Ǚ�f���u�/����q%B�DS��T�#�}A�&g��Q�Wj�އ������j�j�����&}�'BS�7�E� (��J��yfgӯ�Ih���k���z�Ui�-��mڢ��tj�퐟D��\�S����,���q�,0��؜�<,ͪ7��>O�I.�#�ɮ1��ٝ���8k��A`��i ��<��5���v���>��|��/P�/�w0l=j�}�#�*?<��+C�h����3'�C��%�G4y�X�bW��U�0���AM7�qņ�c�9�o���q����"��׽F7������ݳ�W/��(J�#� v����)�S7ir��u�$,��k��4�G�·�f�����P��z᱉I��Z;Q0d��EVJj���-��^������ �f�������˹��ª?pS��>[+c_	�/�)_�%�>�#��������n���s��*P��R�����އ��ќ�#�� ����l����8�����1ȥXE��8���$��F�����L�ws0�,��o���yl=o7y|9��+��c��X�Y�~�u"����A�e����T��EJ�M!y��hݽb�1��Ϯ�b�TRGaZ�W�%�t�����gx9ls�7flڳ�k��y��ŝf�̪�C���6�0E���Q�Z�$3���	��a��k���;�]{�MG�A��ݒ	�1a��He����=z"J*-�X�6�{^���P�Ui\�5!�uz���Q�s���ν�)�h�{��i�U<��}g��^|>eY�?0-( H�y��ظQ֚�A�����-��+Ƴ-a}���qmR�� {�=0
V��_�m��{貙��v�h�ngGM�Db�a�_K@�4����u/�6���_����U�A�$�As�j��T�<H��q�$�4� r�0׺����z�K����o+�(a&�L#��Q(,����@`G�� �/tQ{{����PH���J����9Wy
��' �` �Is�M�{���~�e�X\�9�j�6G��iWHޠ�� J�S{�⊗*N�Y�����H�N���OT0�j0q�?�d�h��H�;g�N!�}���5S�G�Z��c�e�`AM��l�?iE&���Xʜ��<��X��\�s3 lJ�3���ޕ|��S���ta�J���5s��_��g���l�5Y��U?ݱXg�L�p
`v]���d�5�?�=#*�"��n��KVÒ)��,���-�E�6�Q����|v�<:0�y�誉m��uݑ��G5��s� �r��L;��5����
�J���IAm��t�L��Qe�p�P��g����Ţ�B+$��Й��O��Z=dlK � `��J]��OrԵ
��%?^����+�'��6`����xD@j�N������6`<�,�)���
~�H?o���,M���@�(8aF7��QSk��z�^z���gJי�O�ي���5�c�I-�b�_�k���m)��&�o27���x�$�^X{�tjR�:�������T���-�����d�� ���3���P���M�f�As2N�"��hV���_��pn��+�Jo/Z������$/!��#(�zi�#�$��8�G,�AC�*ӈ#�}2���Ĉ�5��a}�zL>��H]<�.F:�:�Y�֑�ѷ�Pk������&ͻw�s�TZN��p�����-�uW�	UC�j^�Ⱥh�M�遴��ȒQ���G��;�����7���$U�_�K�&�y����dqj9J�gsHy#��Dkox?_�]�Gc
�d����aWZZ��9�X*X͖禸� ��~c���{P^��KV�P��Jǋ��}��9�ɴ����a�x68G���3Y�#�D�[����l��a~wg�3.̈́��qz��cg�+�Qk�������3%�B��a��� ��EW����6c� ��r�Z����y�y�1->=`�ӵ_&�s12�=�%�_1A�#?�)���p�m�L�B@pp3�p��E�Ka�b�D��̕�0�$��c�K���\�.t1�E�����m�"v}�`�<���z��zQ4r�B�����I�5){�֫q����^	�,l(��&��*Z��������:��ԗ�sz�Fr�,�6�~�\[����%�I����������4+�˵�t�$�>ZВ] ���7����e�5����{h���M��:����Io�WvC��_��i��1�%&`��O=g�Rȡ.k!�{��E�!�?j�c�J�LVF��j�|~��\����39
c�oեXˍ��f]�BDoI�W�������
�,���N�8<<8?{��iA!`�W=�_�pT��.����眛���82�p��vI.�v�HB�8��<ZoϹuz[��r4Ű�P�5��|j]�&<���z3~��X�}9�[寵it���32�!3����DB5�B��D���j��
��HT�߶l��Ю&a�x���AQ,|��A���$�!W���!0��b��肷pe�H�*�u�M�h��wLҟ�Ą�߃��i8�^�>�O����Y3��^�Հ��G;u,%����6��>j4d�E�c��+ȇSӯ�������A����1Ţ�=!�MK��<e�ﶆ� $UK4(�v�K�O�25|
��z��Z�ԩw�ۤ�痃������)V�E���a
��䌷���u=gF������v����6ka�E/�BXW�s.)O�K�������k�?��g~��t�=�{�qw��L_���&R�S����W�u�΄ef0�Ժ��p�ހ�C�S������ �t�38[s��\��{/��^��+����L�7��f���X�|HΌ�>S��?�Ŭy�'�%���U򷞢l�Z�.�ǽ�/.�$��~�7�a�k��@V;�r�hW���S�d�n��nn
	�Ġ�x��I����<�f��� �W��C�
RR#�ۭ"�����O2�GY�s�
�_�*w����/L��Z��&ɘ��=�N�3Rm1L6��W����96�� Bƭ񾲀=���m�Ka;6�Ź˛�fa�H޶�~a��-r���54>�����F3�Y�O�@���g����Q]cۇ٭ۦ&u�H.᷒�WǟFT��?���{�7Πp�o��_s�m�.7x&5P�n#����q#�&�Z�|�R�C'����7�.�則��?�F�TZ��g_(o���)t�/����0�wx��P�[˘���[�J���GM�����w׸��ȳ��o��J6�]�v7Ǐ�S����h�lE��Іs��S�^��_ޙ!9�0?���*^���V��PG�/�;*����a0[~zP�~����?_�S�؟Ɯ�6��a�ڛvb�IU���[�m#h�(�D��;b���#0�4�GB�\�[d���aݺ�lA��ō��oE�K>l�~7_~��f
��e��������G�u8!��ٍڴ1���ă���3GŻ��I�����M#Zڂx��e�'�d��k� ��ue�l������Y^�N �C6����H��G.[�1@sT`����2����D��K�������ĠX�b����&�|�~4$��r�ia訓?{\��l��),�"�Ȇ1�CO��2y�l�O�L�\02�I�װ����+��@4ޞ9��A�i���{bc.|�%�7J��f16]�� f�ʀ�?&�]˵��I��$ϓ��g E=WI~�$�&��aXs(�J\��x���F!�~��C�zkv	��������O�oSmR��<Tl�IG�ݲ��_!�Z"��9%/��o�4y�⩴�_�	'Cy�ק����c��wmlE �0|f4"�'�;�%��������űl��Y:U�}�sfX;垲�y��qq�FACJ�_3�l��~(���?:�@�4�4��T1�+6rc����po�jJTQ� ���n�K,7v���[���=zl-�Ə?�0K�j�H��>���n����}93:&L�G�������brj޵��>�M�^���:N:/<��ǖ�#�~�gX
�&	�5�*qti���GY�%~��+���g�p������9���Nn�}�ޗ�/�2��rg6Oq�_C ̺��</�G�%��-�{�'�XraR�J�W��D��b��k]��E-
HQ��f�8p��Uz�'wt����o��a��0E,Ȭ�� ?��s���ւc~	xp$ֲ�쵘2����Vz�U4�1�[����	U�O�����T^~4 ��r���f�J��~@Zنf]TZ����x�&.�8(ǅ����pʚ[�
��F�]DK����7jv/;-ظ�������#h�U�R�? d$�x�$�����>�G��j�}��Fе-�$��;̝��	+�'&�[��H 6(�i��{a(����.�W�D�����i[�}�n����wn��2m�k+�2ٍ���^:v��'���k�C���3�x@Rc�}Ҟ��Z;�L��G3��J��Oh���y���f�8ƾ���:|���/+��[pG�[�Of��?C�ǧ�pţu�w�����,�&�����_X	˔0�{�=m��e�C־p��[�C��C��ow�;XpH�7����LZ��MZ���F9���R1S�n5=x?km�}�&PTD�:l���No8���"|�
��żn��ĺ�������P�f�����By?r����v��B�GhY�lio�(J�(�Kzߦ�8�"m#`�WM$��:>uKs~\F�_P�W۵�	'�[�3�0����ň�v,�iǇ��A��c>O���,L�ҏF��Q%u�_�m1�o�Qb��W���i�ITq�-Ù�4�(P���Fo�~aX�4����!���$l����"O|��E�ɲ���7z�Q'"`��O)M�􄩊��E�Ps�Q��k��4 �f�=_�G�Y?�2?
i��6<�A����%$��qaT�r�����_������Y�3%@2@�sCԯ���.u�֢�^�|@I�Gv���~�ms��qz�5- $�(�ן#� jfA"�%B�ٟZ�G��'��k%�Z&�fM�|������%pn+.�f�>�斑1!��؆-�T�ܶ<2*���֭�׏F;�v�(��-5��x� ����\��S9���W�ݯo��;4�T�d�11AMz�YJ���S7�v��}�%��?�fa�I�Fݚ�]��E#���\���ȡl���p����ǚc?����~��/X��R61��'�h1��Z�~T}�.պ>��O�f�|2d�x�[ҍ1���fO�`�6�c�/���'��RR/̾d)VZu!�j��� �h�V��X��R�ʍr���8L���(Եr��=����~+��f�S�fɬˮA�oiaRE�8~�K%�9���l�VpjT�12�w/b��ed�S�E����p{�2�?�{�|Yğ^���`.�ׁ�V%f��;r����GH9,xyLYiN�M[5��%��_[�Q��E�a�~rEv6�koi(��\��쇝os���.&yE�Mg��3���8��.T�ơ���]�:�%י�)!
kz� w ���Ҟ�J$atu����E��W�����S�jK�.M��������������Q$8www.��ww'�C�;!�Ӹ�C���ws�}�8��h�w�%s�Y{U��E���[ϴ�	�E4��z ����!�|ݰw��]��)��Z�;Fm���gk:(+L���"�g�	��h8zQ�Ы���(d�����B �#&���wf&���ؿ�3T�X>,���U�7��Wf�y���g[�r^����"�8�2��7��)�d����3.IAx��������q�f��[��z��! ��+?�Z�e~l��\^9��~&�#ؘ"�M�R޳P�eM�^��H��_��8�G�t)�?�~02�p����������\˸Z�Q]~
A"�wyl���ڀ�w���W!����J�
��O��[���[.��A�%�� ���-�.�KV1�>��*�q��&��}�T�}`�^r�b��jચ�E��)(˵ �S����t�c����mM#�Ob���������pXa���>��G�|�+���@���<�g�k=���Z)�ۿ�N
��`��
㥙j��
����'IXENL<U�v��w���=#���)�D*��	�"e7{?;�ߪY�kN�FW���[��e�F%�F�r.��Zl1s�m�r�P�e�I��d2��2�P]�w�?�GF.FK��9L�?wZy|{<duo۲8�@�qY���oL�F\4���#q��D�[���S���su�?2��\���IKfl��~���gO-Ǹ��{��Y��r7�h�|po�|]|�U��FZMg�7����S�(sJ���IF�x�_�ixn����@˘��Z�|_��߈��B�s�[�ZP�4K�3�s�I����}��'���
����|�WBO�N1I����}�"�]�
}�^�L��o
u�҉W��.w2o��|�X"���<���?P@eս|Tf��o��?_��͕�ğd�A#��b�9Ѹ)e���J5gZu���V�aqp� A븈��=�ĳ��3�S�{+9Z\k���e~�������w{���� p_hޏ���3a� �M;�Ѐҁ8���R����p��|jŘ���զͻ����gau!�=����~�q�>�ى_����f/ʹ�U�ߴT��yba.��e��������dc���G�P����G�?jAg\x����,��,
W~�c��C��P��^����D�U�m�����_�/��:y�_�Qەw3"�n*�������Bv;�-
��(б��9̠��L��? {�0}v>�֡�xw��sȟ����m�ODO�dL�vkQ�lhk��b\Y��=��}]�~�o�9�I�1P�| �3�*��;���4�/��h��k6���o|Er��q�4����i�.����ۨ͏-����sI���D5�:U	���G͏�I\2�Er�`ե���<�f^�o}�oBmK|�e76=�&w�	={]C7|� ��̲����+9ҧ��(���q��V���@��;[:���E�4�i�A�K_0X��O>��3�QxvjZ��k��F�=�w��(�����y'8=	f�6���!���J�|�����g���'����q��K�k0"l0:Â/�����ʤ.��ֹO�,F)r��{�ւTs���K>���cUf�,�Z~9��r��j@�q@�%�K�I<�'= ��=�΂R����d��{~ �z����x+$l֑Ч�;����[�	mP�z�|#�&G�8k��������U�/�y����w�60���S��L�%�:����l��7ю-+�z�	2u�����}ib�Ы��[��k��k�$᳼��^
�{N+�hM�"�PQ|г��d�h�(^z乢^�������t��m<�f^�Ug�i9 �=�$��p��:'�h���'D��>W#V�ì��:�!��h��i� ǈ(�k���
K+|ki���ꆴ�[�dɵ����`�<��������E%�}��፳|�mS�LP(;��r�G��5�����ԁ]d�	+����ЖȰl��ul���Y\���N��P��383�n���B��>)s)C�fj����ص�������]v���h��S�iW�A�7���]�V�a��qooPZǬJߡ���1�@�/t��o		��ӏZ��x��g�L{����'�I�'͡���LO��&��(5�%����'�4�f�*��)a�	r��,�D��O�0% �|\�)+\��>������.IwhZ�y�5�61B����?5Ɏ�,���w�K]�������.�]��"W�N����~������)X_pܹ��a�]��R�Y����vý����e�Tˆ�q�EˬÏ�	6�K�5�?�5���{�l)?	5�����4��b�e��S�
{e�z�Ri��c����������r����k,���VM�����Zv1���*��U�V�π�z�k{���K����ӍX��֤+$�Ԍ�H�/�Ͷ{���S��F:�~c��A���F����Zt[O�)���tN��Xa��zO��͖�Aaz�R�W����GG8��x�U\J^��s���NR�}�3�'�8����Q��t�W��/�[�|b�.�j���}��!� (Z<˶q���� ^'צ���i��A�$���4��-Û�I��|�.VBS{ԫ̴��;V�} �\�(NX������^�2�RR5x)�� ��J��ﯪv˥d�v��?Y|�y�n���~�#����
)�x=%E�5J7���E3�_6Vmus!�]�_c�}Xz��^Ds��!kF��8�� d�U6��������G<=�WD5�������������)�Թ�}gnF�!m?հ�����Xl�-�١w.�y��Z����v_��mm���B��������jNY���IԵ]'&]	[��N�?B4��1y��t�=f.˽#b�c��K�m����ϝF#�� ����2P�*t'22f���Eƀ33�K������\ ٟ[��Wn}&�}.bc��C���ԏ�T��5�r�V�'g���HK4�`r�iN���H �n:�4)J��Kh�*[`�g��~c�=�T���S�qc���I�N��ϗ�⮋(Ǯ#*��$������V����k/�i�B�J0��Dn$l֑t�7�z�8�T�/Q����P�ty˔�9R�nw���;Ɏ����3�z�3~�KY�,?�ht�X��Ϸ_��8m��� �I�Tu��'E��ޯ_r�q��e�%^���{����ܶB�3ު�CK�H�+���Ι�#�����H��_��i(����S�PN��E������8T��r=����2�1�=�Y9dA�ϙ�s'��5���D���s`'nL˚f71��Hs�2L䋓'�7��b��A+7C��6�H0�ʵ��pT����k��ll�S�������2ä!s����,���%cD @?XJaV�������T���8��_�lM��C��z	.� ����3�ۍ����F���ī�D���(w�'�d���V�+�]��V{M6��b�^�E���.0��j�Xn03Vq:9Q�-�_�3��`8������9��@�<0$Hc:6�,~o_ D���
�K?6���u��vb�(~܇���t�rq��'�x%���Ov_�x\��,|�B�Թ��f�9]��oUG�e��=�A���|8���a�I��}^���~Ռ����@ɵ�F�#�]蚝�� ����-sG#͉.��`}��@� �;��j��yZz������P����� �N���r�5� a���<
���і_�=k����8[W�/���8�ia��Be,�}+���[�'�����h�ԗ=݉�(���I�����GR5�dg@q��,���I���E�4��:V���5!���Vv��I#��Z�x�r�Wp3���o�CV֨��[����$��oN��Uu�013M~b�����ÎT>�o�C���h���)+R������A4�w,���x@p�W�tzK#��l�Z�tW��4�Ա���Xq-���*
wg3"�H[6k:�2@�0���?
��$���Vf�t�����]"_���o/=R��Gz6G�^jW7����\��}E1D6��X��M�x%r� 뜾��$� �aQHk��\�	�
JX�L�ԟ~]'�|������1��9�ۥ�9;�X'�?�D��Jɡķ�G�%ac���EςwIt̩1�$�XC�^K�r]?[tY/\�k�� ��
�ܞ����lU�Ϲ��2ٿ�Pķ�E�ݖ�<%�����Db���!!Ǣ���v�Kb�j=��>��#�&̃�ҦInǝI�����8���D@d ��nY�9n7�+�DWר� E�M��a���a�������6��?0���t[_l�3L���(����w-/�%�>���/;����g.���%�����1�$b��q��"Rq��e0�'��<A�#�'z�[��Ղ�3�zS4�{y�Aq�}?.
`�o��[d�r2I�p�<P���5�a-��ɑ��5�;y�d�����Ҳ���	Zɔ�>�*�"�-����*��B���B�S�6gϕ^	P�#�	���,l`bS4S��$@����u� �&ͿEJ��� �.&x��0uqD�өT�����<���+�<̨�e��qol|��3�	��9�S�5}2(�@��k��M>s�s�K�s���%�#\q*��CqdY٠^i�Gn��/+<�O����5Z��N��P���wL���x�8WR��Q喹��_���<��ݖL!O�h�0����G.6m�����q�&��f)5Xm:`�f�^4m�m8��(�>H3=u@��߫�����9��~	�P��A�:���ī� R�1ɿ�?�륆os;iyf��� gԆP��e�ןL>Xn�u��� !�gd��}�C�D�0��]�x�p9
�GG�D7��|L��
SVSlTS#\���=��S��3��\>�_��xNR ؞z8`��
������=�*yѐ>I>Vy�ݸv��"��I���%N'����<�)�a���V�����s�!��������S�?Jkh����'qN�w��g���+�A�B�����+�#�5��5��`��;_w�|`a�	7�>��>�WHbˑ��a���~N��R�
�����1>&�����ԇ�������9�w���|Ԥ=?�Z�;e�rޠ�|��οw�$P����	�G17}'��gF�]�w���$a60i?���<Kz��9��nKz��}3�~�az/fO�w�� �+�!�������@��&�UJ @4n�&y�28 ��
�8�AҎqQ�?S��(ٽ(����/��>���`�uf�-��a��P�Ɔǡ �{ S8È.�<��7������{E�D�F��P�(p������u=�3��� ��o�;C��Bƽ�:A�$1�kT��iW@��~h[8T��\���T�[Ea�F�Ռ�<��32��sٸ"��(�6����M\2�w�N4�����J,)lظ ß���oL��ċ���_ȱ���z?�V�5_� �)���z�y'� ����'���N�/z��H���啅.3DZbPX�'�h�u�:�mi�mDmP� '�7%7 S��VB�
J�C��db'9yʾKG�:+�P�@g`�2�Gg��Ht�Z~��a���ƙH4C#I��7�Ԉ� ��:��cqU�q���W=�4�ϑ����l��[����� @�xS��F���||;r_ݦ׭��"��j�Ze}�>$��àd�gW*Kw�}yG#�I�/R? ��X��#�nMQ���*M�md�`H*͖!v��O��vM���DK�M�\�㸜/��9��!?�����\M��89B�2#�ŸZei�(��w��i|�,C)|t��f�X��P+\ZR��0?�|L%��[#�_�tv)
� ��Cy&�]���5�GX|t��7M���V�F��������
DX��vP:����3^�_���:Q9 �����0c�݇�׾ofDfX��>�&5�vo�ٽr�r\�&���_��x]��F}�ٗ���?F50��w�i��K�I�a���<�Y���I?��4���1���V6+2�`��]�̾̅�x)����,�3�3 ?�Ml��n�;d>���hP��0yT�! ���|�'�r����ڡ�Dɢ>\���=��;�O#�0jT�&��xb�
����f4ko]�EiXH&QN)�e|(���&Z1BC,'�!Y_�;��Z�4���y4G����/pD���`�oE���D&���ҡv�g�a��S��C���V�k~Ϳ�|0nt(��:��0���'��"�p�7d�oM9";B��Dm�pZ�4������4�2b��KuT"���Y���V:%<u��b�Hìc&M�<�g-s��I������x������I�a�Nn 姇Z<��X�/O"�1�ee�~9�<�m�S�:e�6�8{����װsqOɏJ"��7��
����jk��n �D���f��?(x>Os�̚f��0��l�)ǹ��|�j��/�Oz {���=��i���pj�@�#��@�b=�A����L��S��r3ǯ4��ƅ4��JaQ�<�_�a�
���!B�L���� �F{�k[���v}rNy%M&���`na�Y�d���,N���9896RV�穎��W�*� �P)ο!��������`������_[���&�U�#TT�NʂWk�|޿�3�G�Ow��b�w��;~L�i�97�7�#���3�s�Ғ�B3�n��b�������> 脦r�ˢǙ�qoLzZF�<=�Oģ��Oo�_�6v���4TJ���u�0������?�1-0�������OđE�9g�9��Z ����
��Aޒ$X���o�j	.39[-WP8>H�Ң�P�݌�ޗB���7�*w\�\����4�N����يY�m��B�/ �/{�b��p�~��.�����v��h�S�u�͢�Xҋ�N���ňLEe;��.R����HGIbu��'�@LKd֣3ѫG��=ʼ��۶l�I�F� cK"ECo��ӹY)���߱����Q[?�5� �p��c���d� �0 �y���7�3��y!qc�ɀ-������%9�s�E
CJ@@%7\n��X"�6�3@�Aw�8�88��)��O������ �E*������93���iY��3��2"|6i��Axh�p�>w8皳�ܰ��W2$�]L�0�m7��Q�96\q�Eʢ!㾳m~���V�\��%�K��8.��լw@/��c�:*Ϊ�P+��K	M��eE�H9!�!��A��d���wc.}����x�Db=������q�w�eM��8�W�.+nw�����#�Y-[�:�����ħ�Η��"�|�M�'B�Q!�|���e�T�]�y��]��i]�����(�Cil��(������c�OI���i�mI�Y2��@V��L�R���wK���Z߸=wzH�9��b�G~^y�\f�O;�e�����u�*ع�b=��;C�,�#k؂�pM�n�� �'�������$���ʉ��۞q�b�P�n��Ж�ox�2{�a�C0�F���f�X+�$��2��}�)�4�!�C�XL8tR��G@1ius����J�M����'(H4���!�m 	'c|��7��y����S�lS"yJr�`>�H;�Zy`;y���J�E��)������@Ѿ�:98�kV��_?�����V����fn"z.�HTfA�*�}���ß+*a���v�V�d`Ca�C�Y�m���SnjM3�,�m��tw��h7����վ�3[��:e����Ի���  �c��~"y����[\(�2*�Mo���{e�&<mM�2s���l��9�����d�����DKQS1���FxE��?�׆�;�����zs�ֈFcG:�{isݱ�?G�$���.QQ�<�� 9)��O�#��ݜ��@,��Dc��V-�E��~E⚞?��H�P[�³��17�$b�|�35c�|��/Q@�Tw�p��#����䎾��?(�����D���Ey���T��h7����Ƙ�RoH��i��3���'��P���G;�����d}�Ea�f^�S[ڽm-I�����v
�ebbxѾ�:?�@}���~tSq���]�͵7�k�yvC�)���L80�X�%fV�s���T.!Z_lQ T�� �pU�US&�p1`�w�S�g���`ѫ�TV�q�6��C��9��;A]N`�D�u�26�������ol����Uh�(\P��Pn�-X���cRk�I�v3��=8&0l�P>��kg���F\�IH�o��y�ǀ�y�����-��*ϩ}f�}.���L|�~� 	_��[�d�C�`˸����~@M%���D����uA0�h�2 ��i)����ЍY���B�zf�m�s<�v����ĆkM%�M��Xz�kdM�_�b
�fQ/�t�N��j������ƇiUX޾��
=�6��G����E�*� ��џ�RR_T/��)��0n�ZF�0�ōVc}��ԭ�u�n��`(qv�����hZ��d�:?=�O��1?��>�Mw�0�?���yb���	<��Jx��0�J/g��3�x� �#�[��C�!�x�X�ǋ����.�g��lW��`����rb;��G��vZ{;��g������|ƒ�x����+3ǃ��L���<M:vaxM|�Q�_�lcv������/T���n(�&���Zd��������F��CN��|%@�e*xp<�Y��{�3�������s��S��d$j�Va�[�-ɿ�4koM���{ �H-?���D��)%x�z$% u��UA�A'�-��Iћ"+��A�Кa92pF�m����u���!�=W�<�t��G�*�PyR<j�]Ì��6]g��2jZvCoE��1ϫn�Aj���[i����n�����V����'A5��T?  ��Fq�{9w|F�_�o��3P��D���y��y��~9L����ۆ������D�W�"�_B��5_EO�W�f��$k3�w��n /��?"�kh��,�?�.�����}�N�<Î��\��/��-	��@�y\S)��Xr'����<��צ�מ~\mk�L����MȡI������#�e����#���z�:3�v�$����b���; ��m�I��! �)������ ���s�`f?L��$�'����k�"���+��_FvI�*[�ϟ�y��غ�Y7���?�ps��j�\� t���u:7h�e�a����:$�؏^�A�c ��+���*!�0⻕ܣs�uc���A3�g#��J�R�p�b��)��Ȝ���⸘/ڍ�7z3Ʋ�"�����WEY��.IC)��s>�:L�,h�&��A��o��KJ\��5�v{9�-}s{�4L�t�9�t�uw���}�r���U���baE+�lM8����.Í�3��`4P�۩=� ���}���ב�T�{��]=t=�+��)��p�o���&P��#�@�v�� �������*���>	�fA{���2��ZW��,Gn)��@N��w�������\Ƈ>"t�Q58����'%y\:ڂ�����	���s��) kw����Ix���+LZYa�����m�6$ͥ�̫�~%�YѲ�i03�T�J�/c��Hs��;�K?if�]�9JS�Iq�Wr|vI$�o?��Vƾ�_�������a�'yQ9��H�y���;/w�*�߇Mb��Y�ǖ�-���a\䣺���H��ϗb��9��=�|����������K]Ag�6<��́�;�}e����F�Zr��+~:������ʌG��瓰����(�r�ݸ����珢�l�V=��N��ڃ5�֤�(5V�Ӿ+�5QW��%4b�G[o���7�|�m��cӽ�~�ِ;���;Ru~q������D��K�1u�ձ���R�h9�m7�1����>K#1�]��o]�-Z�{�kʄ9J'�q�3i���FϤ^��|�Znj�K_�Ώ��a����M�5�ʏ���^����#��&=��M[�7}�U��M��K
��-pi�I+k;���֣�@0��6��э8+i^��[���]r����=V&g��`�*��qLjG�o����O�Pp��zd^�qn�n�.q+�5�!l�P2�=���#;�,��-r�B4*��D$wU��׮��-��S{y+�������wP�LU�i��v�1��:�l�AX<U��'׺w	�E��W$���s�����
@�;���,�w�!d$�l�>�Jp���C;3�Z �|��#~��{��'y��L�;�0�P����:�'y�#����g�-J��}q��XA_�7�Op���J0Z�p1)J��z�i�2u�
Y��ś�j����/j��uh�Y�X��'��R�FR�51�'>��m,#s:��d5��gu�/B��S�Lg�h��@ؾ
������P.�L��h{#y\=�'f9N��.���w&UG' V'
�?��n\5�طӧ������!ϗݓ�N�AR��n��UW�<���o���e��q?�}
 ������y�jB&����Ϧw���|�~^^�*�d����Wq���$�)��+��U��LOB��zk�ٴ���uۖ-���i9K��H��\�����6�
���4<��G܏/L�W3�c���PX�]��e�мOu�=K��-Φ��l �i�xn�O��A҅�l��ѱ���V_�qMK?Wf��TY��?ڎaԶ�M���% �
ȉ�����V����sG�n+����]��F��Nhr:���0�5�քh> .����QG
���:�>��l�[ZS�|���O�,�A+�������R?Q�4\Gꝑ�C�jy���Q;W��� �0��+R6��n�����95��{��򭑀|6�bC4�w�O/E7d����|ïN�r�P&�{{GsT��rMB����&��������5z���\ve���F�@1�yڞ`���f��"?@����<�fr�ϗN�9��㗷���X!�`���4� ǌZ�7��Ѧ�,�I�v���s�	����U	�D����H��T�e��P���a'U�I����׳�3=�i)���0��H�鲛��5���fx��ٗ�@��_��,@���#; SE+��E���	9�'���4�7��w�ɲ���
>����L�e�� ����ͼD7��������x)"�6�d�w��Lj����� �Z�*��{^K>w4!�G�|Eb��Qz��
J�/k���:�`/&���(G��;��8V(?��3oG6���?�-�+Oh#�u�އ�$a��p]as^�y�P3�\� �!�ı�3_��si�%���п���r�]��AꙠ����xv�V=�O�Fp�" �l7kxj�Ũ��h�>���`����y��ў�#���.�֌�c�PQ�>�9h9�ϺC�u*¯œ�L-T��R
n�}"Zc�^���8F���v�V��uos����zj������9��`���kp�i/7h�5pH��ɶa�eȍv�kӱ@�n��ze�0 V���� ��������F^YN*\�3VJO#<R�)js��j�]	Z�����C�bY���ˡ������]L�"���p�lm7Ǎi5��Q�Eڿ�1���m�V��Z�dͺ4f��d��P��4�Je�I�%����P��|3��D��Z�����$�a��Dӵ|�!����ƭ����hwR�F`v�fH6X�;�C9�3��<�y��h��6D���Z� L�k���ZR3�<��_�Ǩ5���\���KH�����a-cĭ�ѫ�"EME����}:��	a�1��[ˈ|�Ty؁�잎n����龧�x,�>x�g��[�ڎ�F:�~
�~�����ܺ�;��xR��mK g���4�n=냉�t�=�v���/h��e�Sr7hskyu����c2!�`6�L#��o�m7������,��2�=,4�}#��"�ؖ��[5��1&��Ih�E*��qGM��N���	�����)bKŌxO͇7�S^z����J�P>L�Z{sF����S5k�V��R=g�6>M޹�؎������ť�w����VT��ߗ�<�u����DQo�2��i7�:�� T��M I!�}>�0�v��zi.b�O!���bؑ���"`��O�q7�'������}	��ۗ5���dK.�h���D#(��� �M�!�<�$�ȅ{�m�����W��N�I�lv�<�ryQ}Ř}�/��Yho2o�<�^����Z��� ���F�w�6��	u����ώ�d���8��~{'����&7�E�����m�uȜ�ZY4��3ܼ�@OU	��ݱ�BE�B[U���_��ϼn-D��֎�_6?�pE��ܓ�a�� />6�(��Y`�2�T�Tϫ��Q��Mbyr˚�����x>G���Җ�߾w'��<�}����#�L�<eH��R��+^9_� f�o͇3���Y/^/&�����[_�}��IM.ƅ�4ț)!LU�s�!���i@�:�Z$X�°~�|7r�C�:9�x��BU���XƟ)v�\,ߓ�5�.�/���QK���A��#��3�K��7�]0
��Lt]�U�BsIr�k�ѺU�#��N%�^bð|�4D.t	19��7��vU4��D �����������6�a�8�t�Z�L�;,wΑ5d����M;��?�Ȁ�0�
��2��9R�/^]��W;�����ֹ
�wR��X��Li�y^�� >�þ��� i��*��l�7��N]�H�r�O�m#�	�^�YV�ē��5����&F��2�� q����.K�Q�����m�w/� {��?����U�M��_��<����*� �2`��������g��ȆŇQ�v~�4�#vF�m��~��X&q����;�:�I㌕+\�ҽ���9f���9�x@~���[�m囄�x��H�j���,H��Ҵz<�{x�s�������&��"��7F6�C�{�7�gS��n9ZX]����*M����܃�a
7�{��*c�80(�nD�ܑ�<��,0g�$��a ¨��Q`��ՑO���7z��*o����G�X���&��[cǙyq|��Z��x�ET��i�.�Hk#���A����^,�IQy��/�N��h��޽�]�73��GV�Q>��ګR&k�}��H���`F���	/�HG����TI���C֏���s��ٺ��������FTAϛg^���D��ees���e��I����a�����٤��a��V%#�n�N�ɧÑ:f��NA��?��fV/���� ��Gc�����@o`K��!h���H@ �ʨ�I�k��I�M���i�o�(�3A~�~��&Z�5����S�6e����Q!s3i��b�������qXXѼJ�~��k �����U���\x��^�klv�N���$P�K�����x")�g�v|{�z{A8t���Lz����b��P�3$/$�����翆���j���	��z�)0y�*��j=��p{o.u�c6T�"���#.\]3;���@B�������v�-��op�%�e@vJ�$H��{}rvg��WE�x�%�V��&ai{��`
����+���S�F��ꓚ��p�[�-��}�2@�������8S��cAY��m�(~�;�g���{��!�k:31�C�4!�|P��L�kF��́$�h��r:��y���%�����x�)
E'�"��!:&_�i��gy�% pF�k)�l�H'�C`:jҋW�P�S�O 3�#��	~1��󤛴;�i�>\��C�$�`/�-������n�L_�e��ӻ��1�{��[=��t��Ô����<Jko�O��av{e\���NF���-8�4|>�u"�+����V͛b��������S��0}}������eN,l��ī[6�4���I�D����� 8 �������~N���5x�R�D���R
=�el�#dM),�;��:zo$�A����i��P�<s�n�ؘ��x�"�}3�撁�(N�h�e>��b�cv�S_�|*K����:�����T~S=�s���M+�6:萂�+Ʒ� _ׅ�̥�Q,7�X��f���s�"F�gh1���ч?Stf+f�_;��CJ΅0;��|�}>̀��+� Ġ���#[�=�uQ��R���RG��ֹ2��Z��&S����QHf����w�Js���f��y#�~u3b���<�|�m��>(�rd���=P�T訰%��|�9<�!�p�i�_���c��13;�l��Hq����[�<6p���c�5���/�=���ָ�懪"�|��kMfoc+1I��z��2����g}o����⥰�Wn[sW���O���Bʕ�ۘ1��n�)nMu�i�cK�r?��[�Q�,k��&TD̎G�^�5�^$�\xL�b��+(R,
�MH�G	'��<�^����s���O�noA/uB�8#���V��B_J��#�hD�zM�[@�hL_w���^�$6hj�n�Ѧ��ҏz{Ŵ���=��F�2_���Z֔gUC�o�2�� �)�*��'4�^�$]tn�`p����(�~�֏W�KZw{#oڹ>�}G¡�,ϕ,���k��.��q]4PZ�}���xsLL�+�F��2�iM��E�]�&K�e�h�c��ǑV-z�x�
jgiZ�Y��N{���{a�t ���O�V?�po�O��&N��'��K�K�������L[n���9c��fRXH�ɛYmyd!o�U���j4SI�S�U���
��N4�c����Z�̈�^��Ұ����F�0��p�|Nķ2�^����m(��ALkD��!�L���$��k.���-Ey6����a�3��>��Uc­���9bВƹQ&������N���F��0W�Gu6>����{u��j���Rk6&��^~�@��5��D� ��KO�T�u�u�G��R������n�֬��u�@��h�}�(��v!��F�u��a�l'~��2B;u���y� ͉�cO����n4,�r{�a����ͼ�cʕke��.���} �� s�y��z*�b�ǨX�)���ڐc0)���O{�8�v�^(�vk�Ā�Ll�ꦗ���`AՋ�س<�ǫl	a�D,kr�VZ��
�jt�&L�k�,�酿��4�/��}g&����ȯy�y��$d<��N�67�&@9�y�u+���U��n�k�<O<�r>h����6���vۨ��5�j�^�/ئ"��,ԭl�/���y�<�
��:�d���A�r�c�rM$��@��a�L@x�[�YO��Y/	ol�w
rZ�狩��r;P�G���|Jv�&�.D����9XX�?���C}dS���ڶ;�Z�����: �"H��b�,��}ڞ�HQ^Hz���$��0�
"~&�ǆֲ���h�撋I!�4����Ͳڏ'#.�c�7���ס�	�}�t�>{E%��s�Sx�:���
���@�����B�VJ�����4����Xr ��W���<
��^���fU�t{���o!�H�#�>3}�f�%�����*�E�/?�1�Ez�ůa{�Ïe2 >�5��� {�����#Uu�U���y,Ϧ����m
@���x��'�6�@��8:��8���4!#�79�'��m���"�s׿t\�ⱛ�5���\ �g -���:�Po1���g�pA�&���'��+Aާ>bb��).�b�yB]n�K5W�\El������򗺪OZG�հ0a1�<��,6U��h��&m��w��S�J!�m� QZfVO��z��z�'�z� ��W��*/�1p:w��l��@���%޶���/�{�v����[ǜ�����T`����E�G�J����0�Ԅ�N\���2�_Kh��-?:�8VQ����.�z|�s��L��.�t��P_�f��vBB~��P���e2��w�:����.R��R,2���H�i1gY��^��-ȗ�����nϽ{?�����������k^��sI���U�Sӆd�eq�^��Ro]o�-�_��>�����L��O��y��Y��%S��48�|���|�<[��韗F���[>jǙnlӮ���b����Lhَc�t3�U�sQ�j$n�љD� "kS���˥��$eA��ٺ��*%�Ld���*�H|P�}�5[�7�\�O���	r���[��^��~�a� ���Vb�}�@�nzV[��"�?�"�∜���&vܵ�6�m�n7��t�����rl�bA��w=d'Df�k��7�H�pq"Ւ䛫���
�J8Wy��E���\��FvI*��͹�R;5���k:^� �P&x��� �����1֬b���H�w����~��o '�7�����|O�3��L�x�����o���AG���$̥��K��>� �Ջ��@P�yA����/ו�\�d9��8.��9�f�ణ������4���^R����*�ʂ����%ִ̑jË������,.{)�/[Jv���n&�'P�42}��ZN�ZUָ�tzET89q�xFȍ@�5�Ȳ���v�@�hd�V�^~�����a��?^L'���WUsxg48�Z�ַ3Wl��y�� :���Lw�,���?�{G�&~䁴��M�����,��O��4[4�a�/@�2#��tK��C��΢�a�7�aa���Z�^	�4�"l�����G�YF��5[ww��.�ݝ��$8���]�Cp�`���=��s��[�_�Y�f��T�~v�陙��O,�Yt�=��)',�ط	�)%Ca����ͺǕ���8ܜ�Mj�R9m5s���_��h�~����-��m�yV�D�;���?���`����Ay�)����t�$�[�m|'���}����/���J��5��0�٥�x����dܯD�z�
:�O���̟�:}���}��XL%����dސ����q8���/� �?�c%�U��	���cH�X٫yE���#�Ͻj��O��K�#�GV�'��J�.%2Bu�W�E6YD#�"R`�r��h�gOFV�c��C
�6H��|J��N�[�+����� �v���C��D3nsyuc���^6�3z�7T�|���r#B��	�=
Fp`3E �H��Lc'f��d�h������H�+�H��p~���ܺ�6��z�T�I_({T�p�+W���;s&6u��.����aC����o�CWx�+��(��0PP/=@�n�yo:�n�}�|��[E��S��R,R��m�	��g|@��t&��ͧM7>'D� J����f�tj09���sf��Y�Y��m�ќ�����>��w�����R��@	]�=�컽���J�&2��Ŏ�� ����V�����
?:_��h��L9��QxC֠���9s�3u�������Ì#E�*b����@3�3��aˍ��E8T=w��Qa??����`=h��ʛ_g�̈a})�)x�D�<z�`��ӝ�y�	��n�ϳk�n�&錓Q?��Ԥ�B�  =��:bI�b��9R߲�����d�5ڻ��/��]m~�?��:�2~�r�֓�Gӵ���LHW��T�]_�L�pwr4矙���'n+�wogqn�Gd�MQ�#�B��N]B�4��gp7Zw]��0��<���A!��;Z��=�λe�}��˛����m+@/.8�Ƨ�����Z�b�&e�>q~
��ҭ���OW��4��,��?�RW=Ԇ��gtA1#�-#ێq�q�IC� ���d�b�.���1ccR���$������2r���뗞򧑽��(�-%"�\Mk�,۱����	Rܩ���$P�hk���7F	�0k��#c�ՠ0�@��^L��X>�[8<�8'�컊�d�A��0�2à����p��#wU�@��E���`�#��\h0�=8�n�!�"��8(F��Ť�Y�p������X�<'�T�JT4�$Kn�>_�(=��wO�3�Cۛ�֒�^5۴�M�Q��Ъ��92k � >ɠ�D���9�?wI�����$��'-���1糠��N�S��3����K�v�&4k�X�R�T/؜�7hPb�8N�콃����*8�d}�P�Q᮶ �U^�|����ޚvɩw�E��K��ov	��Ʌ��`X��aX�S���+��>Y�8����,�O�o�B%��l'���8��������Q�=�n�_�m�eNڛ���͆���f�3o��$��⦌��8�7OMDB���7%�bz���x���]m^)��Q��<�q��A&�B�f����	
S�q�?Hf�G��I�3 � ��1b��9����s:���;�
��u�X$@aeb���2[	$*@�3x�S�O唇��h��1�{fd�����
.�'��G�n9%Ss�Ê��� 2Wu�B�䘏��/��caUt#���U����.���f�Ŀ9mҎn_�Rě1�b�u�t�C��N�fcF+w�[z��I�^��,|X!s��Ɯd��9:�7&ݯg���c���o�j�����R6˼I�r?�ɨ&-)�i��ęۂ�x>�(�,zz\�����0���	tۓ6��c�&y4ޯ�Җ�^,�D�?�"��X$L�F���v�,�P�Bo�7��Z$���P&%t���J	t��T?������|���a`wo� 1��3����MMB|�>�������(?Ƅ�AӇ��7��?�~���\��*�SK����>��X��˥�}���g$ui�����+�h��D�{���ccd��p�i�O�8��|�D�.��x�~�.⇲&�W��k�7��{eS���%�a8|_��3��������'��	, ��ԭ��5�dչQ6���G9�$�8��`�A'��W�w[�Jp����c��ϣ�_r:�E��$Y�_kLN{�J��"��Q^L��z��V� ��nN����CCȿ���;d��k�/�T&O|��k��h��E���m&�V<����ݻ���;g�!@3���dQE`<p����aR�?*�e���W�@�	���?���y�868�i()_>�m1Y��r�?�O�O\T��6tfStm�Q�����1UЭ�X��8��/�GB���撖��������Z2��:���ſ��[GƦ�"�e�	~.3��@B�_�߅$�gW��=vs�d�}������.k�Q�V<�h��k�w&b-p�3��N�"�f��%{�вV?���4T(��|�c�a�����X�����U7�G �Pj'��Ll�q����D���������K����$k�(�gh}��3��%:�3��zӚ��ր���m�F���xy�]�p^��Mu�{,��ͤFˇ�QP�����2��{�ѧ,lŌޛ�dĮ��8w�iC����/�Gc��&4Z���,��ˢ's����*EBEN]?)��� ��'e�R3o�oT�bc�	OͶ-*(^��ƿ��ȧ{��{1�΁��+~���`��
Y����F������[��i~��d�!y��f��_h *r<��� ��7mg�S�@@�G֦�nr�b��������� ��v���|�|��;#Lzq=+�眡'�CPI[Ԡ��3�i�V
�J�_h%P#�g�c��OT&0)���~��8��%yp�l� 8�J���D��$uZY"��j���e����r��u����"C�?'^�*��_}C]ͧ�`
������ � f�[���	����a@����+�r�	n9W�6[>e��*�w�τI-}�̄v����l���7	Rj�p�i�bEX#T�4���a��!����H=H�V��31Zc�=���b�������8t_���B�%��Zaj}��lb���!{B�IF`R.��dhH�Y]e�jH0��.o�t}M�+��BS�yi�����j_�1�B�*3eR�l����E{�j����J����E�dV:o$��sO��ы�C��uy�Tm�ɩز�B�C�h
���r";)ь�Q��͟��V��l�w�<���F��$H�l���9�H���i��S��πL�p��ԫղ��pG�����F�f�P1sg`���G��d���E�nl��S�M@�a3B�g��_�O�6T#�'<v����R{}�ac��{,�r�	$r�둈S/�3� ��a@�3Ki��Az)�~'�� �G�TUF?g��uy�8�*o��D-�����Z|�uT��|���K-�l�����c�P���JgǖğT������m$��n-�Wqd���2$�l⻋����R�j�Z	�;]�S���Pe�fϵ�� Q��6|���0<ot����3��;g$嗫�����%-��t18bв��,L�|Cx�p�Җ%�QϘ��,�j<s��C0A�V����
c��t/}��ӣ�8�� �x�������zc�3X+��!Z�a�|]�ކ0z/�N�)wh�ﺧ���q��چ�u`訧E�?�;��u��>��AFV~\��a�L�i&�S���f���|��f}�7K����ˣX�{A�v�3��q&�]��Gq�~A�taذ+آ*V��9��h��A����5� ZV�]�r��_�;;�`�2d���RqJzpc
���d��������kr>nƔ���w�7T�QԸ3ӇT%ɂ+h��@rvMn���LKsJ�c���ݣ����ᒼ���H4KN`gL~G5���5ǻ�u%cz��Ι���u����ͅ�
9��6J�_�S�[!'����qx�i���8ڻ����{����B���DDL1&�Nx�fv�Bt��n�d4�C�Q��Cwux~`��b�m�BV6��9	���(Q��sq�{u-��w�Z�}q~�g�<P>
��2��Tc��^��g2��P�69Y�И�.�E��o �#�0���R��R� �Kbk�@	Q�y��nz�Xo�T������YK�o�۴@&�͌`!�%MC�鰥l���S�W"aJ��E��n���iՖ��6sƋ}�AGv��#�
	FPq	;"pZ}a��[/��c��"�V?���eC%ؗ�<*�����PG���OsSNM�Cq#�����O�7�>R�p=3@��t��x���[�6�
��
�Q�2����s[�Yi���t��Y'o5�p2ryM
�q��Y��Q,�@�161L��6��:�trx�Qç�1�6[o�l���8$���9�"qd��"Pkr���]\y�IV�ʅ�u]Q(�#��ͫ���� z9gV!�/�D)��9|�4 �'��⳩�_K�k�������~�����~�B�{?�v��8#0EsӞ^:�t���!_� ��<Ls<Q�!�0��:J���K���ӧ$tS֞ �D���k���1��v��,���`���M��r+�A�X��n	���^�gkcV��R��ގ~�U��J
�u�JU��D�_ޗ�;\Y1�M��vQ7�ޙo�vm�;漿z��>��~��+;���D�݌��W��얗��Ө���ўy�?6�܌��,`�����.����jN��!��>8+T_�gK� �	oޏ�����^#�Rj��%@��N��W������j��D�=��*���c�6j�f~�P��`�6�Іk�rϞ���6:�-��[	���G�����">&� ~:e.�j�� �F�5r/d�E�����}��ZH�3h�[��<3�� �-��d9�6G�o3\�} ��m��K*yb�Po�CT�Ԗ �J��\'�XI,%�]U:$u���4�2�bqS�&3�k�����Z���^�����8����y��\���L�3��*��W����#�:���IBw|d�{��
�/�1Br�]QCrH��9��y��
O�L?��ôa7�fc4΄��>��r������G&{u�︐��r1/��0��$��{5�B��9`A����W#78ma%9�ו�}�3�qrv(8�{{�WI��G��ֆm-M��ƹ��;�����d���l����nR�D�<�5�5�0Z�A*/ԅʿ��:R��D�7��ՅC��$�*Yo����E�
�B���}��$Ml�R+�w��# ��$0g[!��ɚ�P�a�����EBº(QH��Xl0aMD9]�	Hۃ�Q_�	L� ���Tv��EhY��C�,������p������ �F&B���Y9L�̬檘UՕSy���;��:a�I�Gx�+��zs����؁�E^=cW1�@=��'�W�v�{��q�ο�LD�ľ����}�⦛]z�t�/�PЗ�y��$"���1�O? �f��ް��W��/0w"�5bGR��k���@����������@�p4�l��iꢚ �f�I���*e�9�z�*�Sב�	��<a�&��	��E�����`P;�}��|J!
�L�Ά���jީ��aف�b�ϵ��p��-i��:�䥱�z۫�2bk8b��o�IV�sD��n��qp3�pT�9��%O�`;:ڽ\��n�
Aݜ�����Y��/hdz��&�݌�e����~�Ri����d�e�I��٬a �<ϷH�Ǫ8�t���j���S`7�E���I6ԲoE������0*7cS#�J��~�	ꤰ��^�x* |2!�Y�iڞ��<�����1��p�Z�B�|*q(�?ӊ<�\��&�E�up�:�PAɈ��M�r�����.�y|�PܥR�s}��+�D�1NY6"���
I������n��s��+�N�
o�g��²D�	[�V��EdN���z����e%!��@�Ó����0?sJw��2���ף9�����`�O_p<�[�����-�cM%W�N'^�G�����Pf��>S�lbA�}�]�^�G���I'%�9�
���m�j���>\��dFVo�Z,FC�����-"K�h��.|��|	zD�ן_���"0���Ő7�dZT����1����~U��ax�z{*�Z����튮�
�x8�F�\�����,�> d�吇���Kh7W��
W������C�5����\���ON�/�:+�gq�}M��^�AĞn��Z�~�\_'�d�*�h��F��'r7�Ȥ~��LGp�z|ɯ@DPs���(��0�L�X��i���e#�)�c:�.���ՃNz�`&=J��[��R�s�ۅ��`)^L�/r�a�u����T��@P~5�H'LFV��#��$�`�!3� ��v��xw�")OV"݄�;E�r�W=0�ϵ�(|�nc&a�t8�ߔ���3�6&�|I������M�.�fL��b��fk	��/�-�������ja<���4��TV:$�����m��}{�"	�"Y�8����o��A�Od��@�~���^��w��_S��^��t�����1H���F�3֡U,���ɥ%�ҏ�M�h·���n>{%�ƴ@A��t�ۛg�/�˭��C�����]V�ڡ���j�CgG�U�Z�*�M
�>Bt�n�[��S�
�f2g	�Km����ODI��A�@u�N���옿TM�s�[v��d:(jI�+��\o�T��۵Z�rt
;�ɷ����E?�Ԋ���<�����;g��V�AqY�V�}tKH Cmd��*�V��e�F3������ `����мÐ�A�D��o�I%�ijp@�r_ȋ.���M���ޮ��<q�1��4F��۱||����gJ�õ�A���#��/'���}p쫢Q��h�<��Q]nc1����c�d�	)����ڵ!?̃����'<d�~Q8�'�6��ܛWp���\��c@"���׏�t �c,����KϿ#�m&ׯ1�z��e8t��P����%�����޲��r��srܛ�"�ڣr[6.[1�+��`�GЕ��X�����	;����fEd��W�銒��x/<r;9m<�k�z�K��S����u=jyJE&K�(���67���6˺}Z��7��S$\=o�n'����M����UЃސ]�řVeݔ<��W��8Myq#���ՊH������5�vɋ�o�	X<b�x�ުji�q���0�ef&���gB۱���;�$�����ӄdy�-a�d}��!���jAI��b٨�������5�K�K��`PLQhr�5,��utz����>�0����`�I����	�Y�K%K{ف�Ǔ�������d�57��;t����(X���$܆�}�3/g��!�F|���#о�T�@s3�5� �d���)�)���)�w�&�)vdE_�f��^L�ZH0ȯ�޸�m�ϪD������wU;��� ������#Хb�:.v�)�<Ŗ�tP;���Q@jҩ/׆Qrg�b%J�%<�W/]-N�t��B��d|�G����MWzq�2�'�(�˄����޳>z���R����}�ٗ��"m�"*����1Ȑ񊞹�p%;��-Acd���(Օ�����5����d1h����z��
�&x�F[�Hu�u�%Đ�܆̞�l�x��~�XK�kL]~�4em=��D[RM�M>�)��椡<Y߶O�F��E�N]x�*�w�OYeGw�u��j�h�xn�M�_�w+c�\t�~�G�9^����}�]DSJ{�~%q�Pa 	I���p/�>I�kXd7`�������|w�%c;8�4������[ʟ��2��ݦN3">�j�QE����L1����3`/ng����#Jk 57�!vT�!i�2���7�l��w��ȣ���ׯ@c�aQ�f�|�2)�KY�Nv�M�@VEJ��U[�hMt��C�ڣ[J6�v�o�.��4w���p�7O ��!���:ǖ"\I,��	����3�f�EԢ� ��;#�)��8��! �>�/>�.��2Y�ߨ(y/�P9����"�J
�02BNv��M��냶p�����)�W�c�Ǔ��ఇH{m7��x#_��̨|5�{�[�;r����q�gg�L#l�ڷ�Ț���v����N�*�O@�)td���b�l"�z��cH�ɹ�5T�圝���6 �g� ����"$Q�h���鼍������Υd(���Io�B!{ғo�4d��Z0�d]�,l�05]�-����� �C��L�c�^!K �C]�Z���l��i��Z3!�9�dCW�R�xJ�5S��%�&�?���Ѯ�w��ᔷ�G�a��������A+	��K5��فl�,�-%kR�����p}lz�:
�D�]�3<V��+z}:gC���5�e�á��żǽ�5Ej�4����>W���)v6�G�A5��B�j�E,��>���U�n�-�%��e�sN6C�e3#n�#��dhf�� ���1���{Z�����[Gi���s��k
����{F�<n
�,ֶ�$-ωۤQR~�F{P���í�R�ŘX�_���Ҋ~�̽U�RCN��7��*K;f]��J�����I�	��0fhi.��j�IV/dP�|g�i��	��M֭wo���u?Wu�`%�*^j�$ȩ:ʕ�'�3F��q�%��E�ցk�;6�)�$�b'd쑚��l�F�`f!v�_�ڒ7sOǡ�z%�a�SuO�]#�ˑ�����xj0�(I��$�zF��o|�?��܇����tU��.V�|�n���������^��5y��گf�v@]�{z�rv�^!B���N�(ؽ�=�<
�����,���\��T���`�SU^Mܠ��헴�a8���~d5��q��ֽ�,)��v^��~�p�'�}öЛ��'�w���z�zg��yr+�CYO-&M��F;~�=�2ߑD!d���/��/�rP�c� �9 �G��B�4Fg�N��$/D�Xd�Т{�~I�H��ܚ4���0�������|h�֒:���;��:���y^w���c5�ce�LC���Rk�Z��ο�O�E,�yN�v^����2z���+�G(X!<��,�o���,�u(���3VAh�>� ����/��f���؃��_�c}Dz���FP2қp�S�I}:2�n�s{x;��9�l9RpZ��� ,)>P�_�\��d7��>'K��ߤ��|{9�FDNW&�I���-r�A�*���ܮ��]Ǯ�
��ĵ����KM��eܴ��։�y��Dދ�K�������3�4�Ҥg�f�̊I����!���]9GN����"]�[��I�������/|���5�7P#t��J����5��RV�:�⎘�}C�����.7n(~[��n�&��ٱ��;�,��Y�Ε��������t�M�,��:����%��^j
W!��K��@�Yb��+~�,w��BV��7��\N��-b�Y�1�HI�(e|�d���PN/�����%���=i-@�Ԯ�,Y�����ˉxp�/|~z�<��$�Z#�>&qr���h����\��4oc* ��k�`	T_D���Gd1϶_�ŋ֎��!DG'��E/��1�O�HT�t�L�q�o��A�O�~�u٠��Rz�L��*Zx;�G�����l2�+Oz�����	`�h�m/�(��=��7�RGe��ě����sr�4WlC� ��x
����ɩ������@C?w���*�s���W/�#�����.�	x���KaK�L�t��|l���u��`%)��0H�V�v���
rE9����C�T8qZ���-Ґ�'��gE�@���;�9�qR�I��1����-�K�	ބ�&�����d��|���O���H�Z�V�b׃*��K�r8�I��9�) |h�+���+s�nw����^L�^ٔB)o�$�E��1��\���%ƃ��ƙ;�?�6>�;�/}I�	c��Hv攀rIF��!���m�������겵�5
��w"k�@KT-�Lc�35t2���4�/3���6��[W��>K�l��C3�����ƫ;�-� ��0�������D�9��5��0ڭγ��"�]`��c��X�,9��.��n6t�~u/� 0Ʈ�g����%.\����_K�t����u	=%�Y�,��h;��6I�������^$.�&�{�B7�����뫳V@gI>tg���ұ&)C:_o�&C_ٌ��q�߈�������K�q��۔,�ڦEa,F��� �d+��Hd���-G��!i?|m��g��֣sb;dǵ/ݮ�}�H��3�vF��7��Z��>n��$��J�Y�'�UR���t�f��8Ӑ�`����߁�(�ܗ�`�����Wn$Z�y�V\Gv�
®ίڻ&�zv�v��f�V�jT�>6;=�殠n�2���Q����Q6H��!��:���
���/8ST���~�LB����>����Ѝ�έ�����|X���k'u�����`96 <���t����\����P��kӋ��e����1K�V�"	�I���<׬���a!5�=Z�q������z�bؾ����昵M,Jܫ������O�-�t��\���*�S^ɲ�-��jh��{ٸ��s�p=�ۭ��'n�mn����v��o�>��D/��F�����U۴��y#�b#��1���v�|��a7�@CS�/�s�-��Ի�d�1ߓ��� �MX;�!��5���^Q�f���1���g(l0M"�5���h!a�������T��_���̖���zJ\Ga�؜�c��vܐYm�Jd���񴼲œ�䧶'�C����I�g��ē�\�I�j�ؿS�f�vb*��3�i;���V�qʔK�y��e;�=�I��D9"A�m�Is��z���ޏ�
�1ɼ�i0؎Ő�:��K�s��7�ن�vB3js�$�'�n%�3|#7�_�b�&뫣��^n�]�L-�Jt(�3�q���D�N�������vN��j_>v�<.�*��O�.
m
�����tu�aE���C�5��]hI��mR2%�~O��+�f����^;e�����d�}	X3=J��>�@4��?��O���U}}�X�s`~��K¶Y�r5���@@��H����u�����V��_G֧����\�2"�HD�5�g_QB�Cyu}@P���T��wf��%a�~&��<�B ������.�����5�S����mN)���D:6�^s�r����B��H��}I۸+L��K®FR~�N��9�d�cxמ�Bn���![�ʀ,�\���*���ߵ��/�|��A�� <��y�@ǫׁ
ג}���<����ӝ2T�~���_�`��GH�6!�n4|��.�D��L�k���epQݹEP�����mx�r*��D�w�Y��o���t�J�^4��S�GK�lQ(iE.a�M�=5zi���w��	��"_����i%#c�sC����j�M��1_o�|?g�w�l�N�5C�K�36_�=,�2��]�&�y���Ďl���z.�P�	O�jWϸ��(���I����2 �Z�h�Žř5����@�$�}�k�m�]�X7�3��"#E�BOQ�r`�� ����i�� ;f(5�����3����_H�c>�K�\�|��������,$=��]G<�M� �oOy��P9�j9.k�_�]'��&�R|�}�T������oDH���XT���a��E� Hs�d�6��$.[�h�T�i݉��z.��%Ug �������:ۚpWF�r���fz�I�����f����g7�6k�����턾�zQ��*Q���i!5#�a�)p��C��bo�ݔq�����@�m(i�z��[��RHܜ�bc�������&��&4��>�Q�ѱ�^��Ӊ�>�� �M�A�5��(�ym]
5'8O[���jG��l�s����y��8}�x�ʒ�����EM���`�Rg��r�%�2B S^�7G9 ס*�>o���h;�<�mT�Y�9H�J�a�����M+�(�T���l����A�"��9���x��j� 8I�WX!*��r�.хl\7;�o�+����N�Ѯ� ��ـ�*p�@�(�6�UG4%��A?ܶ�����׼Y ���HȄ	x�M�RV���mJ��& �X�R��J\��?��wR}Q����a��	HI�W{QB�l�ُ��Y����{�Q�bm��r����N����9b�lɺ�8Klb�>�*���H  �����8��.t0'��bg_�p9��㩢*n�����un��WݚT���k��jΆ������K�d��T��Q�.Y*�����{Q����Y�tY��īH�m��M�[�:�@�M�(Iș����]�"xP��m��o涶�{Tt�x����<V�F?�#@����{�
Ŵ��^v�4��h��U��\��Ӯ��Ż�D;�����95s�}yHW��������V*�NEpI�~��sI�D:v��$��	�0�/۱7D?�^B؎�f^�U/�q�Ѵ�����.�Z�۟yy~��3�P�[( ����j�O���Ҟ ����!� ���Բ����,'���	C���"�
9��y�>��N=<l��W�1���2����M`���X�U��xJ�&1j"2'�����`�K5�:uB1��Pʤ����ިr�P�1A�V�Y:�_��͘0�$���P��;$�B~���s�-牖� C�Y�m�G�f����b����J�MF�� �R��':LH�L��}��	T�M�fb���
B*�/�;)�uBk�f���Y� ����FP��^׿�ϥ�0�D����%����?�X�:�4N�0]��#ks�3�����ц�=��n\��d7��A�#���/��\���s|�Y.x�~��̀�3~;ߑ��8qW�U-V���Q
ȟ08R�lVbߕ�:���y��U�eGP�b��?ږ@�6k���t6{O^"��B�x`d�.ݽ��M�xw�k,|jj
1@��9V|��;�i���u%����bi�b"=�x^�^j����"	ۈ�0_$U��]������+R�k��ˑ6�z~��c�(��I:s�����t�5nPX`��4m��<�j�1�� �3���=�Z7$ԕ?�c#�y����q���I8�{�kxmė�b�M���7�6��,uOK�����j����剩�u�C���O�*&8��4SC�Um�yu.p��T6<����d���0�0��X6�H"�q�7�ϮFDx
��)�^�5�0��?[4=^A�?�
�X��5zٜD ѽH�찚����`�o�~#)��L?HNn��I��*Q�L�n�5��&
�ۈZ��ٷa)���K�/�dG��9����.�fh~S�R:�b]*Y1%CO�e�F©��	$�>(-��.�Ɵ$����=���E(R]�0{0~������&��.Xp��vO�б=%���!��b��
�cz.3n�TU$j�?���׊j��`�ī�`;�ʯؼVW�ي�*U"-�0,yaW�� K_f�ސWWN���Xzj%��(�p�E�a���C��u-�t�˗��o+�Y}�+�(�q�Ic/�lP�t�q�3�urL=� )n�
;.ǀ�3���ˁ�C��µ���&��
�_���|��d�@^,���s� \���#E;��ۧ����;�0)��/{���I�>��`�jՎe7�ڻ}�ާ����8�x��T�ɴ�N��5`۳�^��d^�O��'���O���/A�����/�j������%�0����@��!!�A3� �������C[tZ�I�OmD)@����oeQ����P��VSFHQ��{�6�A^
�<D��Y7"��es`�J�ř���V,��������?����U���m�,��O�ίV���u�~<��">�dz\~���]g����TG�l��(�����~��:�p����\`�#�͟\�����AI����:)����47�R�7%U
����زc�̸�ڨݐͷ!�!�,ם�ۣ#��2Y4M4��ж��gmn �v���5��_ޜ	fց��Źhd-��[��W�{�Ku�hn�^x��Y�A.�U������]���I~�ƭ��������������"���ܝ��J�)2%�AZ�e�5[j��Gx�ΡڇD�GD��p'j�s"��}� �������6s^P� �r��@�Ҁt�ф�3؟�`:_ŀ�d�QZE�2��S(�{n��h��>���q�	:���P�'(��^���z̵�.7�:?2��������}`yv�G|�Q����ZH�,�W١W�؜�1����I�>�_Ļ6gCW��� "u��@E��Z�n�~�z�v�5�T�����}s����f��;��M��WpSh*2�/�Z������?m8u
���0|M�5�,/��I��V��A�g����=�,�.�:��O4k�ja3d)�]Y����0F&���#9�,��z¾�<h�3N��A���Q�`���/��$kx���_�t�SG����:R8
t�ڏ}S�meЀ��^#��ZmY���md�?��p�2_t9󾉶;r';Up8��8<��24H[�����z��A���E�:��>����
��]]K�RvQ�%���&�ѧX�a�8{9p+^zZ%�զCs�s|�����^!���e�v%�~o�T,�!2TL���U=����|�w�Y�nR�\�)��Frh�J�2?��ࡑ����#2�M���Ѷ��}��즻��0$aW�� 6Xc3�rtI�X���y������������%��Ǌ&2n�~�,8�� *ޜk�B��후��s���3�n�LL�̽U��=�ZZ���J����\CD���z ��l�q��R��Ǔou��s��W�eڹ�F�b4���y����`�{7�#q2����#O�^pa�dQ��r�nQ*�3T��
�a�%�8)2�q݊�c��Hhxr~�脷��ُ��j��f�!X�:��]�n�RГ��(���>r,c�-J�@1�o���B�0V]�P(U1���h"�H4-��{m\(�'���P6@`I�	B��L��@�`,2=ek
3��ܾ�=�)�e�jZ�� ���z�	���|���� 	,��I�Uq�f���L�ܩ�bi�I�2�X���ufژt���*�P횯V��K����sǙn�W���� q�	���p�
��	����W���Q����(���%���cKy�?qy��-B���'�йs�<M�t��6��˪��^��o��~��'�l�"P r�n��,*~�G)��v��m\z��n���YH�g�t1���1�e#�}qE��E`�5����9�b_�x*�^���X3��q`F͒�(Je0��^~u ^6ä��m�CQ� ˻����-�����H��ϧ9'��/�@CdEA
Q�0@��ЄlqŦA�@�A���t�B ���Ѐ���+#���twb��r$����Hpn{�E��w��������k�' "zM��h@���n�dz�%D���ey"�p"PK�����Ɖ��{(��R���K��@j��sښ���<�Mo�L����h|���e 28Kqh+��:6�V
�ʖ��YVj�2�	�[ٗ�rr
4kZ{�A��7�����y�콽�C 2M7�=�8�b]7;���V�ʅ�%��P����Kg��9/�XT��"\�m�-Y�]Q�W�mu7ε�J'�0��e�	�YƙF���җ�n6!�[]y��U%��0Q��7I?dWo�#���v3�T�,wK��ش���T����1�c0�uV��<���n��kZiC+T�dG�v�#�TFWG���&H;L���*J��R�e��ppCt?c�!h��W��ɗ1Cf����(X��@�uY㊙�5�MY���5��={i|>���e*Q�Q;n���F_�立%2�~������U�%���H�E���i�5|�?p��9��K�K�ߔ����0j�x>��p�b�BQ9�c��3����u�I����2��Ks��hŇ!*����W���1D��U�)b ���),��o�r���XZ�5^�Y�SL:����<Z�����-2n�*%q��jw��Ĉ;��s�2z���Kiܡ/����֧��pB��(����gD2�l�w�k�q�����F9E�jE�B�tʿ��*��[��#�ƛ�X�f�%MV��ɶ����P�
M�I`\:�.2o�����	��'٦.9�<�u6&\<��#���� �N���l�o��4��á����E�Yi҈��F�i��,�,Y]�>׆n�ςgF7Nr�Ԝѿ-��di'�<��U>�)^�B��ʞA(L�rȮg�p�AGYKlCS� �����տ�׼h���N�f����Yj�N�篲K��8 �S�݆0c�悢���K�?I����t[V/68{.X��K�/ۢ����|8ސ�e��Y�dQ�%w�<�1{f�k��=c�ѵ��nF��n�z꙳R�?�]yO{�T=D J���H" H�m{�����l� ����-â�ڶ�ABA�A��n����A���n���$�a��a��=���~�����xg��X�8�c?�}�k��R�퍣�rľu��t����U�0�
��{~L)�e�Au��C�ő^�j�?Le��
��e�l�����5�������%�w���U������=^��)���>��_�¶Cnr��G�D%Kq�f�09�����C��r4�C�l���a��ɏ�@��|]X�����)��Y�����m�`���47��5�I���}W!*#�߄�׾�P/��i��b�����	�O���g�4U.wv�l2��Q��NRx����cA��[�X�d�mq��ZlE�!3� $�x��@�:
L�*.�g�������X�&ʷt�Uu"�cj����e�蜅����p5����>����'9��J��*��.�"���{%�+!T����o�>��2[�Oz!��&{���|1�j��2��V� �~�LQ� �П�@r*�������^��h2�W� $#!�~�9E�]��'�$Z��M����J��&eJ��P���Jd�\[�ƨ-r��_-S���@�-[X���w5%��0�����53c��aW<�M�� ����kٲ�ˣ�y��P�Oľ�pW:��n�P֊����7	�A����(|OR��1ЌWW��W���]WVu%zm�n�n^t�i۝�O��gd��H��V�r�vą���I�F�&��X?��Vjf/(?�!�9_���x��g�=q̜�<v1�JԿ���ӭ�&�R����WSz`��J�<,�ӫ{R�.
p���;�H�S��e��cu�!\��#E�	�%^3`���k�唥T�	ÎUrth���uZ��}x�Ɋq�!xS��w��ƪ1�;~�\ʹz0!+\ʈ���8�S�V��X��.�P��]�+˗��#ړr�Z+RAا�S�b��Zm
<=���H:�=7�[�`#��K1�a�`R~\,߰q�P��_����%���� �н� �?��y��f[��rk3�nu/��M�7S�<�V
�x��~Gt���e����F���PX�@���klEub����Mx��	OȬ|\5S�Z�Ux��B�13�`پ$a�FЉ�W�'P�N�W+�Z�<�W˟^�+����Ч
z���J�����L���U�ܘQ�F���1���.9�ؖo�EIG��hd�����t�&�Qu�[�&W��e*����,�-\�DH��P����-�0������j|L��֠��+�_Y5������$7�4 �AD��lj��.~�\��v�6N������fEQ�����Y����u����c\w��'�5M�=�J�j�MZ�3���\�D:�E%���`�@T��v/S1Oqm��B1�:���M��T��߽U(����\��=D2�cOim_��A�0-�c���@�욋�u���(���l��n{B�%�/�����j&��x�B1t`�˭,�L�Aϝ�c!Wa�b\�Z_*�㞥�Na�6-N����Zg;$w&v����������Q���2�RK�*}C{\�@��̽�/��J��e���w�K_�$�X����o=� ��m$�g�w�����{��<���c@��)�ܴ����
��V�-��IOe~w��1o�v�$�˖�[y��[�{Q�8=gZ]���7��v�CGry�1�T����Uəͻ����E�L\(��4}Y��(�>kdk��jl� �J�U��Tk_��x[	�JE���`:Z|�\��J�����	E�4t�Y��E�eh���eл(k��۟䱑��C��n|B�����ݷ���)���*eof��@f��5�i� ����P��X	�Y������> 6Vݜ8sްCr�"� �ѕ�%'�`�Ԓ�x����K�0&�X��}�.i/z��a��C7@�:�	#��Oc%�s2�'$(�]�,z\��~/ʌ�6������5v��}C���r��7'�-����v8�U�[���X�����7b ݈>���)n�6�7�S��v{�c�O���`}��� �����S�ȏ���i��l�7l�(`Uu���)�T:�m�(2�F+	�d;_��ۢ�����V�kW�T8&��q�j��c�nRW���$�5l*m%I�ޗ;�۔���s7=������o�6��$����Ĭ��s�ԹF��ּ�	P��N�"������RtӤi)Ee��o����ьA�tb�@��*�����ʺNE�.�_u aDG?�3�O���n2/���e������2��s�&_�t�C��9��~P?R���'ڍҜ���O�%{����T��5�-M�'�j�4��j�:Gj��`�	���4)��%�����O���+Jn �.x�/F�+ K��XRo����|CD��!��vt���,��W5�����KR"O�nZ��/f\,�����^���SDgVu��z���Z�Ы�����Ę�\�ܿx��	x�T)�)Px����H�K��������
@n+m��[Vk!�p�D|�`�w�@[h���u	 /��?W��B���Ul��d�2�8w�R:H�
�7+��q:�K�� �gm�_�\����K�7e��-[�� e!�����tC���`{~Fǭ�Қ�%E�D#��-w@����[!v��`>�Ӭ�����yM=�W����M�   ��`���I�
�L�M���"�BJO�L_��5�1� ��ӵ��T'���[��#I*�7�:��Vce3�w3�m�m�[� �8?�A���E�x��[��İ\���:s�t_�5����5W!sO�O�o��q/�y�s>9^��=���d(n��M����p$��t�gS�a��3���ZT���8��^�t����U���|J��b^�2�q�*���*���̩G�rd�|[oI��w�Cn���g4 lm��o�{��&�R�P��~�þ�g�:��D��|�E%�ĺ��7Uf0��������g��ŜA��_h�U��e��W�?���z�p��}n��,�wQ�n��/qO�5��ُ�x��A��C!.�ҝ/VMЩs�;��H��ř�T0�jy�����/*�P~r�d X�j�
���b���V-�� +�[�A���m�iQ+�1��$q�g�_=;�KC���w��� 	{;�JjM'6&��q0TZP-��[N�?�5�_�^�e��������=����ei�O=�S��-�����ˇ_D��*�a��T����[{�kU��ٙ���Q4J�rZB_D��}��r���� UD=H���ѢaYD"r��10��|�q��c@I�F)1/�������d%����ɔI�Z�9/6�pبh����4�y���c] �sF揞ž�z���b������~0���0� 	�aL0!B�9��v���1�Ǳ<oG�� �=,/r+��=�Ա+1�q�^���ԃZQ�Գ��\�I�v�Q]��L�Q�\*�[tk��*�ىgt]�ްd��I���Q:~=�T���W�Eg�/E�����/W�Ի}���fq��SD��� 2%�(s���X�)�#����(K��K^�NpU5��ђ~�F����נ���2�v�g��ȍ�l��3^��ZT�2B�XQq���Je7����GIg!�SD�_���ڞ�4,��X<����j7�Ԭ?9�f�����{ Y
�>o�ן�G��!�[�=Hmx�%�%���<�����f�Mf�GA�?���೓���\#�7�ځ��С|�tن��Vt�"ө�=�T���S՛���дI���׼͓:���G���뉴�"�@%pRd�m<tm��{ڙ�&�y�t��٣o�K�9^TTb�4��/���(����i�O8�ߦ|%O�Ej�0E�����gY�3�a�/��� b�/
4�[���;�	��?���Uu����n��x5�G�J<J8E�� �x��핕�	��v���1͑�,f��
�3�E�e� ��G�ܝ)��Gz���=eL�0z	���S�|7���ݲ��������ǻg#@�ȝ���@�ߪP)��aШN�����W��+f���w��Ӫ�Q�����#?�~?)�C�ﻉ@�P��\��9Im���fnn��
vg�`3=��y�գ�����Ǧr�{M?�V�a�;�" �;2^�Pб�+H�������@:M� ���SQ9�)5k�o��s��_��� m���ߞԚ7�m�9T�"x�4D���C�V/K�!PgT�ei�7��I{�i��P���&�Dq`��t|�f_S�/A:�'��`��xq��q�^��+���鰲�"<{��K�rt��ڻ1d�-rm::�t�Nz�?w=8��c�맋�F��D�`�[9=4�OM��!��tR��/� �Z/ͼ�����4y��db���I�BS��M@0���'�ԟ�)2�Y�d�䏫3�'�a|$hT�/=����G���,>���+�%Q���͌�=G
�I�۴(��L�Mu%�n����V�=��<���(�Q�Eu�!`�?[�Ѵ��˻=r;uY�T��gO������8���G�m%[*j��'�%ot���M�6��Ĉ$���8��l�"���M��͉�.	���5���/L��Y�{�)G��9�	 (Q���.�_ɂ���A�@,{p���mP[�\��N�a��~<�}��N���>9�����XDYw�-/g��M��u���6���8�iv��d�ա��pš��
���|b��:d���C��K��I^H�m#֪����9U/ $<�^�i測8���4wh>bh����W�yj�]�3I.ߨ�+sn����O� 2�BTxW9%�*G���?2�	�<W+k����ِ�g����8�t��?��^�����Œ��é?s�8����9��b����RZT
�D$����ϵu�"r%H��P�r9�T���c�J:]���Ǽ��UVƜ�8<��������G���ˎ�{�}��� =�������O�<!��*[�ch�>7��Kx/�uƀ�)	�x&/�P<Dw�ef|�A�z�ȴ��)!G���5�s�2�w�\��"�<w��΄E:���D#�}·��ӡu�2�#����0)�#���p�9g,���KCB\t�SS�\���O,��f�����6b�X��c�;�9lĘD(�1l�,wv����b��v��eZ��^ B�'B|ק,�FĤ��ʨ�ʘ�2ܫ}�ع����3m��#�I�8���,Zh3g݆̈́f��#��2ͺ�t�i��e��I��)ф�
��h�+ �����������,?��|������u�:Km�͂�5P�����g�:��9���~����L-��}��{�{[�k/�S�v���,���m���|�	3^l�r������N���
����힞�@t�l�wT�GG�a�s&��eUL`�^s��oM��µ��b�� ���S��U���oo/R�]�7 7:�ǾJ ��~�!��K�����W֍�<l�jT5Ru\��4�Qw�>>��B��e�2��9��2!<3��<\��M��<V&��&���erhڠ��5�Q�H�ٺ���'M&I�1gGhT�|����g�;ɸ�D�pe�J\���u�"C�jm�A2�O�?ZZ�r��nm�wbڪB2�⣓AaJ���Y��z�&e���A��6�V�#��
���G���Y���L�[۬B�h�TiM�&���ov�٫/̡�*c��ڀ��7�����%���@��r ����k�s�&[P<��R�Ju5��[�.o���'�����N��u.jX_��ߔV$ۓ9�i=G�a5�u��N��0Cy����<��k���櫅���h�8򿯘^`�}'�������Q��wⰱ$�~A�g��C#-���q��?C���X��p����BP�+!O��&���?���sڹ9k7���y��$��pc��#�ñ+�G�;�<����F�>(�}�&t��������	��PGd��ߞ����ߟ4s����i��i��ֳ8��$D)ژ2�ӿ�>u1p~��V��{3ay�������*��������>���Z�o�cjY�����t����˂ǵ֏��y��?ҌSXҜ��@�B|�R����Ь���m8���ܭ�8[����ʿ�z����
�i�i��Xy��L�S%��@���. ���/�������|%?��{I؊>�+��ļ/��79����4)�o(�lN�O��ī))���H��>n�p��clZQ�Q%Iݙ��U�DyT�mE�LLt��iIG��N��De������?���/�x���f{i,��J+յ�?o�i3��:/-��U��s[پz..���[�dZ�(qQ��Ci�<�W��f"`+25�AEMO�r���|����)a���o�3���f�R��1�f�nɮV�d^�����ty� 3AC^j��9�r��w�d�����e�/�9`�O\ο�Җ��eO}�;��[#n���^j�*o��f��0_A/G��4z(���ܞ��I�L��O�󈔧8�&y�0Y�;��j���[x�Ș�./�U��]J8U,�V�8kz�AA��D�
�u��2u���L��~{��V	0! Y���ͪ��<�?�I )ߝtx!�����㥪�N'�lIҲR
+<
�p��3������a׫����������"��H��A�y����J@�pϑڹ�r���Y��֠��Q��\	�_��L�N^Ș[%ʘN���j�}q	��;-I>o�c�h�G=��(�}��^��^�9xV�⢻�^#ĩ*n�6�*�w����h���%�E"/ GO�*WB^��+ݶ��(� �%�y!���K�Eq��qmc�&�61b�>FEߍ���"B��|�u>�v�����S
(��H����H�m�j�Y�L�L�
���0O5��Y2�~�H�*���B9�����\��H���	���3)��uѓ|�U󠲼"ҥ٩�˼����h�r%'��愤�u��T�8:����g�������jI{��	�����a,�b�H�V�>�~�Cv�T��siM�i>Z;汴D�t�Z�S9���~IY�ѝu���D�*�B�����0ӊ�osu��������o�;�\eΌ�R��k����"�|>cK6	vn������2��y��9y�F�{�#2b=u�^���@6�����;�'����'ᐉS���zR�+��w�K��뼏�s�͡q!���tdꇀ�z=ݣ���k��:�ך��/�]��7����e��4���֏j7KFEf�u_��л����­4�*m������U�c)��5KdMX�^���śz��»0���@���ZޟY�/o�Sw�#iGq)�Ǩ��Z�D޶�g�@�7a�C+7vUѤ]��<I��^�������`��C�w�7��v���QV4�zFY���8�2<� ����:�鐚����k���1Y~������N���&��_��ړ��{!s��~k6�7ݐ���F��"4�ҏ:%���aá�`�V�c�R&҅�';�����������Q�m��Մ"ם��V�M��ևS�/�B �9�s�
�bf!I�� 5���U��;� )w�>�^�����tН���)r�hԣ&��	�G�(�c#����Fk���Z��� �9K�Ĳ((�n��LQ�*��.��	��d\?�\��U�(��!I����'�05�_7�)�ᣨo�4'�2��wn��\f���3���׭�/�� ����5{˭��`��a�Brq�k�'[A\֥iߡr���l1���H����UD�#�v��!�%�yJ�Zz�e�n8��h:�T��[����w]�R�M���Mv��Z��_�l���v��������O���֝k�yͺu�U�I���)�D�m�aL	0���wl�M�m�Y�%[�Ճ�+)���	��E��fx�5��n|��iR��j��t��D\Qv��Ez�	�3�U9��^���<e���t�I�A7&��sfXs�'�z����۾�:����a1q��ss���y���~	t#viM-�I)(:P�Фմw{���Q]>�vW]��:�[>/�������C�6CȪr�r.�0�׵���fM�n�d�ǐ� �3�ъ�c�a�yN�����`���fKf�WBx������JٔB[�E��if����(�Y�L�A����~�f��m�Tu����Wd;u��ܕ_?+�Y-��#���2д�\G��(O���uĤ���>����2,6ic�q��$�g<.�T� �tZ� 6P�۳���(*
��`�Z�m�p��UT�^��~��Ɠ�{�7EB$�%b'��IT��:���Q2c�t��Gx��@�s��8x�Nt��x�����p�����=�1>=��ޞ�/'ݻ쒒?G�����2FCfح�ҏo���4{b�(�����;�u\��<G�/�	Y�0��w��4vJ�m����o\����}89c��-d���}5�b��&rM56����^o]\$�Pҥ��s�I[6t]#Z��0��:�=,;��Y?�� (�VX�V6C��>c,jx	�����5��|v�/�TW�U����b+0�b8Z-��]_m�![&��_��Gm�<��T�E;/�x���r���N�9<�g�f���U��%o���������U��"xWI�D�q�w�u��ĺ��,���#Bm���NE����du4e��d�<�\~�02��\N~�`v��RA�=S�P���R ���X$|~�ѝ��dc���S?0�X�U�$�{[q@���!��~ɀ�V��R2O�1��� �?K��XFM�ݱ]����I3O��ff��F.�Bq�KG���J�TTH\̐�g�`$�U��S`�4T���]�m �-���D�P���v	��S�*(���n����B�f�=��Sݥ�x�̯�+�v�sw�&D��
0������,�������� 7��&#�#�S�T�۱���:���q\*�gp}�f+�|���>r���
A|������:u�!�w-��m!�O�ԵvKP���.&����P�D	9s��z'bzʝ�CN�-X�Ѷ8}��'����
�u�*�_��K�<��"g�#���]# '�2\�r=Y<qz��R��i�% �ơEױ�<#cUЅ�x�*���~�5"M�fN����z��j���h�$���M��H6&7Y��I��
W�؇��� ;*�c�|�4��:gy
�d����	�|[�)!v�3 �~2�\����˝8y����b�"��������-gug:�6z� w�Ա����?�rY��HQV���~Q��
f肇�Ȧ���a�ι��0S�s`�KYK��ZR�6�dS<�{OZ����f;j>/HZ����0�O�.kxE?]} �w�;�*��Aj
m�x*����"sܧ,+�:`Q��|�zx2vR(��@�_@%�kb;u˻@���ה�!���|�­K�N���o�8�a>�2��Go�:Y���E��	��L�U�lp
6I$G�h�sk/
��T��|bU�؋8ʓPn;[
a�TĆ�M��V�R�Tb^�ܹ��C`y����ӓFS���W�nN��K&L�J(~H4�m�Ú�5���rʤ��-���^t��IXlV?��I=b�h��M���X��A�;����}Yi�rm�܉���i�1�p�]-�k��iK��~@ar���uk����b������|�e�����|c�q�Z���R�O���fA�J����{K+(F�<Yǯ��5��"6��n"F��f|-͗F�v6��|��Ǹ��/EzU T��ts��O$X�T�A ���Mi�vh�Y�F����XN�6��a��M��7$�)KM|���)��>�M����%!�#���E�+�\��$� rb*���D�ߊ^d:ս׈Lz�'���{ yѶ8i��>�H��.�,	6vV�����w�`"�Ì��k�����8]�F���ͮy���7�ެ�L�v	B���B��ebq댧e�N���J�f���wԣ�b�����7�m�;�n�|a�y��R�;�#:V�f�;j�s�������GM��I���K�gޏ�^��4e��I��Y��B?j��"2�;���!F����{�.>t�;תRT8�T8�r'�B@�[ZX(O����B�g���7��u�QhP���~�h��XsN{��I�� ��KxE�@o�|L�9���tiG_�F �tp�<���[$�:��6�q�ֿ�k Z/{����� h�冄h{cf��eYr)�8إ	f��B�;����x��A���������T=�&�V�f}�$�7���#��;N��ӎ&@�3o��$h���̴>i��j�B�dJ��8죻H�f`.�KP(��<����g�_�U��"��Q���o$��\��Fk����s�h���1�ͭ��o���T����<M�/���C7�&�e�m�?-�o��)�����N������`ͷ_��G{�ȟ���.ɤ�r���CZa�@����{�o$)J*�%��j��~>�[���X��iO�tr�~���o�R���Gx��\�.R��
t�,�C;��v�ѯ7�6��2[љi�	0�ނ�ȐעQ=3D��	�bۖ�~_<��Zqg��R�C����=;��PQ!�h뺩�|��d>3��UP�z��T<�rI���0wCxUC[�S��<�dKo��]��"���fm���%���'V��>Nr�5+�����_Uڗ�zaL��D��-�$���$J�x�/F��,6*Z�?��\~P��2�����LZp�ֱ�'�<_RL���00�7����Y2��!��B���5ǽ%���5
�' � �f�g��1A��c��E���l$�-�mך�VLT��������=�j�<i�9_�3s1� ��a��u�����8�$�-��t4�N�o�BG�$�d�{���T+����\�Ux{�k� ���?�a�p2���s}����ʍK�`��X�Q�����w���ʧ�$����Q��+���b)��a>�P����L��ݫ��W���%	
��(^Fg���o�VÙ[�^?�|gWjK'�) 4}ۦ�<��M7��+5P�Ξ�ld��qm���.t��\�t���cؒ��݄�Z�z���q��ѯqב��]���L�BKx�w	t����*^X�c;[�r�R]���V�̥���O���_ql!�s)6��+��Z�W�Ȼe���C>�uq�W�nso��@��4�I$K	��xZ��8h�b����8
����[��.��m�4����~ש�^�v��y�Dv���i�Ӌ���_ �`L+�H� ����
�TH��;�Q�%`
3>���b�Lz�y�B��|t�8����9���ד�O4����O[{-��"�+^쉭*U�.�R�3%���.�J�?�|�$J�a�s�M����f�cI�� M�w������_�n }��`��7��-5���Se d/�����Z���~�Xjc/��gb5�m��X�
�W+P+*l����*��çF��'>	�`-�I),ɴ��9*6�P��ԥ;"��unv���	��,Y-/��f�M�8�MoI�?h�Ț�j^1�G��.�6o5���~e���'���i���ĥ��7V�;7]��Ф�<2�f�G���;��C.e�ۄK�v�$i��������{O��	2;�s>�?� ���Q!@�5 zpq�K=��ÿ?)z|��W�-T.�ѡ2�ZS=]�b��UpPo���*̐�9Z-Km
�(��{�@߶;�]��9��H�Tv6���)Y����O(��6���p݉+�G����:�߻��7i��h&{щ�D��{XӦԐ�䛓��+�����Zam�lSV�@�����γ�bDB�>�a�7lڬW"�Kg���:���R�vL�����.&R�뢝i��H`)���绍���}�?�s�W�J)�/�lxZi���?Q�*򏢯W���,r�2n~/��]]�����kJ[R�=jA�ѵ)�9��v�L���3���
2�Ih�kƠp
��j޼����p住�4�zl����&=-6�Lϡ�����N�}�q.�E��yM��0�%��&�,�x��4n_=͙����c�-�3Q")��:;���\���JU����q]��m�HOSSQ�����e\���@H� ��Z�M�/a���n2���k�n|���)��A$��ag�X���g�{՝�,�ƪ��?x������H2���A �[�cU[Z��գ_�����F�ă#b���R�	����r�Ҿ�|�Z��;/iZ��e���e4�*���'bЀPb�2����U�����F[Uh�6\֯�>��V�>��Նٛ�h^��X�L`�,z��3$�R�,�ŝ�Hk_�e�B�8p� D�T�����X���� MMf�v�\ECٳ�S����.F�.���@���D2ӱ�e�^��_��ӳ'P��E��t�e?�9�rU��ڨ��a!�����*��-a�3/�}���c�����`,*D"��Vi�q���R�G����� A�썶�����M����jщ9�]Ɍ/��^V�1����zj��-�Z�����[J��ǺAZ�,�����ၦ�)v��,4���Z�̫9�&���[��LHs��N�Vǅ3��T��Rn�����	����",�3�ׂ�|���!!�gS �ُ�i�0������1���:�d�8�ֵ�d]���t,9��=�tU�� ���~3�0��0�'�����g~-�rS��F2L�Rۅ����cP�ί50��j�b�c��C��}`#)��-�~��n؅BpNA�XI�7��c���[ )�X
���U��y�����H��Ӥ���Kѷ	Z�
8�;�^��gZ긣�8_�����V�6pq��' ������u�]0���������k��R6۟�K���гmD*�51�si�R�s�J��z,% �#�|�喹�'�R&A0~Sz��������M��l`�i��-�g�ȶ~���;!_@����*����=k	�T
�n��Sa��XҤ�9����k8w�rR������U�$W��m+�����1��G&�喆����� �Տ��'�j��fKc�CD#�j��
ba��HG�UԔgҪ��Y^U61�=3�[\,��4!1�]�H'ٻB��DZ�Q��]I��R���6�`�OHH�U�;�`/^{��̚�w&�g�|H��<�=:PA�,�H���f�JY���12 ��%�����Ӓ#������HӳeݎX�3�k��u+f�x����������"�Y�v/+Uv�|XH�9}X���y��M�$by=��Z(��*�%g����	3���{ :��~���L�΢YЍ��-�2G�S���6�]�� �G�����<��
�/k�o5�u�v~b��MU�9%;=s�
M܊����E@���z��D�\b���;��[��#N�l�L��/�����[ !��U��!K���y�+�V�k�<��׾�=]��zs��V��?��^s�^`�P�Y�T4�'��b����]|TW�.����Nw(*��'���)+��젥��IS�p�l[��Z��E�jy�|�db�d~#��f��g4"������x^�Z�n�4ی���s�kV����8��?�jAI։��$z-][�䋇�g1|�^Q�z�6���@�����|f�S��|�?@7}_�����~y����l^�ǃ�G�~b�=�!��+��m������&~/{����<��;��G ɥ��b��M���N�S�^��1��X��/��˚��&�'(z	z����m���׫�}���UR�QZ��>��<�'�c�"g��`�黯Ǯ\)�sJn�oB�e��-!k�s��I�Ζa>�R6$r}Ssc�Q�eU��?ڼN~���m�S���2�o/����=rZ�r����~ �a�ލ��-�-Q5_�TJ���c�Ȯ�Z������Z��l�S���x��L���D��Մ���\�O���]؟�|zw,>A�T�6=�.gc����f(	] �����Hv� ��ޤ��J��E��fK�6y�&|�4�q=s�������� Y�m߆*4�2˨�WMS�p�N��/@�h��恴L��e��̿OD�h]\��C�6�|���1Z<��ֽ��mӇ�1�1\l ~�n<���/���~��	*N!�W�v�7����)Z�'݆e���v�e�L#Q�)ߎR�Bj�K��}<`Ӽ'ô�F�4tWTm��m!��o�BK�\Լ�.G4�̂SZ�Ul�2룁"�nR�#��'o�i����e��&D~m�d��uW��K�h�kip.�&Ɋ-D��]EIy��H\hg��b:'Lx�l[uC��<3r�}�y�V[x
�l�~��l�=w���4[ev���ث����UC��R��5�@E+w�@�?$]E�L@��\\%������� 4˦rvq�3��
2Q������Ֆ�8t��!���My� ���8_��`rISC�b���J�mY�+��*j�����Ҿ q�p��a�x�~w�1�yQ�?	�92n��@�M͓#�u�"�����R9�Bw�$�M��_�u��OEҠgg������J0^�4��� �>w�P?w�`:#6?[^��a���՞���k��z0� U��q�1���
����[�Nv>���3RRJ�g������|'�|�R�!�6i׳l���t���.�p%L�/�_�V4W��^��R�ߋ޻~�7eP~��(�9�x�m��;?_O���?��fwl!P���9n�hu�Y�oښ�zC��&�r_�aɵ�3�T����ZD�6=0�(2{�~��XE[:)��6a,���t������Ĳ��R:�U���Wy�۲}�y&>h?n��'�����������>�G�<�����N7�f%!ݓ|N����۪{�#8П(w|��2�4�ivl����;5�����\��u���&�݂�YR��j���>�@'L=�������q{�j	�y��� yz��1�I�we&)^�E��C��a�?��`Z���¢U�6�������gۊviƣ>��Ρ^R����Q���ۀ5�%��n���꡵Ӯ�l�/����%<���!/)��s�:�p���)˚B%A�͚/��wN+,bip�ݻ�tm(f�ͦ���<��e���<w� �:��V��e۹�o�Sщ: :=��Bn�9�8K��C���}������zU|�{Q��4�v[�?����v�f�� nm���VlJ�>�xf�g���8��m'���>@�>������I��D�?o�-M�E"0����f���]Ђ���|�wAX�ϣG����^E����&�vN��3B�ܼ�k��~����y��˄ss�%�/!|�v�@
���8
�m��0v�2.į*�� +�K��F�[�mcj*W5t�%ZO�P[ X�T����Z��d�v���<��. �����"*WWQ-i���8߱+���-�ɚ��Q.��pyh�Mwh�)�UP*�Λ����e��H�fxxF}P���C�nO�v:�-Qv]���1KQ�+Sm2Q�m�������&x�O�0��|�i�͚�pD��8�r����_����5=&��	;g�m,�O.�q��DŔ�C<+�.7�7y���z�fr�qM��Ho�17ߢ9x�i�q�+�:�0���U�L���nM`�P\����mR|k(���&8�ڐ,L����o��}\�}�ߙ��|����v��Yd��9E5�xF��*��^��깳�r�[������ԍ?�;�B�=��:��u��̜V	�k:�Dg�衊�3��BӲ���(�L��n	���~���+�����?ۙuv�3.���=����M	Cо5\��:/8� ����}A;��ӕK6���Wy_+?ESK��IXY������e�>�۲ܛО�k�_�[�Z����ö��Q����,�������}}`��Ӟf���ᡓ�fr'ҡE�	Y�\��֑�i�P��)@	]��L��>[y��휻{Q�7	���W�g�Υ�^AK�~�G��%v � $�-����h��m����P�b��M�N���`9pK9jL�,g�w�{�D��A�`Ezb��2�|aA�jw�*~�v��E��ֆe�)<����B\5�����a
b�nbx>� 4�wH	�ϊ�PZg�����r�|$��
b��H������t���i���z"膂����?������O��R�|��٘��v�� �Z�MUI��&Ԥ��+����{g���3?:=��H�OB�9	�Ƌ7n���[�Ԁ�BVa����������T�0����pڬt�/�sy�ה9`_���I�zK�w���5������*�4 �I�B�xS��:����0�u�J���?�m*�a�Y���&ȧ�����tUz~4LIp���7�����k}U|��Q�����߁�'��W�U��=��UB��o�$^�q��>�܏��c�-XK���`]�N��B�T�ϙ�״nҢ�夳��`՘��7�h4u�2_L����ki�S�>@^����\J���δ|F�����ʋ.'3Ր�	**Z�
�m����vM�����vLdM��7��dF骲ń�R_��G� �G:�@E� �O� �l�����]��I����� �Y�	��P(�=%̐1�|N�2�L프�'��^l�c�8ːw�X������!��:�ͣΎ3�N�G�����X�ѧo��-K�7��a��y�� 䶔��6_��/�h.c5�êh%%�|}ȁ��|���������	�(�_L���F)�������|�#.�G�=���C֙��r{u��E��?�X�o��%l��L^ە�m�ܐ��.����X����?L|TU��EZ@�[���.�i�n��[����t�tww�;W���YK*�;{曙��g^z��[�Qee��./ء�������[��б@?�7��ܮ\�-z���-�s�ښx�/:�/�f�&�3?�"���U�|����9q_�L�z7ű�m�W���Y���Y����#����R�ѷ2kH��ܽ�_8k7�ռ�ʔ|�P����*�q�)��}4Ë�Ɏ��c
�՟ޭ��J���lwō��sOS\�V���9��XT�y��%��)�u�,�^Z�Ը�s�ѥ{D�D�z���<�f%���́���Pߟx��S��{T���z/�[/Lu5fo^u�k�c�G�^Z���o9/�T.i�m������"G�:�5}ůK�fF�Dɥ&���۱f�8�f��/������h�z��W\�H���I���	��P��g�*E?��
��j�X`�rXY�m�t/�XQ����'��cǸ�i�
��ԏT�'a2���)j��1u�Ύ�$h ���U�贵�ƻ���7
�Υ�^$F6'��I�Y��te�W�����@�$���u����^f�>*N���eOn���D߉�����֎/����6��3 ;\�ҧE�k((�ʆ�3�
���D�l�e�s9����3+l ]��p���� ��^ဦ�D)���]�lZ�w~�����yx��V�t�bB�棽�����%�u!^�TO<V_/$����
��M��υ��]�(��z�S�~�|��`�{�C����4[)�]�7�H?$���Y�q>��}�x/�p7���ְ��4���;��Dk4��	
L�T�n-��W;���j*NT�xd7��Z#����k�#	[!�7��L{�~��u�L���q�_��j����I���A%�ުc���\�η���A�4������'˚4$�I��4���R	���C J��l�4���0�ܰ/�90�N|{U���ü@�����ު렞����d���+l���$��Zd��S�;�����!��qM>�wa��c�и�)ԪG��6�u��@r��!���
v�ϑy�K�.|����˓�=dn�Z�U6�i��zy�,p$;+J���#i�WK�<\%)48ǳئ:OU�-� �斱r��sʌ�]i�$�K?\�:YyC*GчEK!��x��ׂ��/���Vs��R���ނV/9�'&t�8�D�喼�H��,��s�V���p�Mb�&�D&3��^r2x���:�*#�{��<�z������>�oR�8��ϕ�TQ��|I,�j��E#�Ҙ���>��I����ބ	s�Q�Fyw�T�H���������b�QҾ��i�ceC5��!P�T����\��;Ώ�b4� ]��o��&ܚ~N��ՈUѯ\�n�N�D��ߓ��8�����Ќb.��^ ��o逰�d�#�_����!?%�q���+�ګ���l^.�6�^+1���>��)�b���ؖ	�5�E�1N��~�y�`��b�:�@�f[4ԓ���T����9�Nh�.�a��J.�'Os.g�����ŧН���@�T�����4Xx�X�x�� ����J�Z��7�%�a�7I���	� \��S9g���A��H�����B��ê�d�|:dbb�'Y��Uy1s(c何Ղ�$}���1b:�Y����J��%#��o.;��a@8�#
QD+�|����ӳm�&�T�"���	�NJ��~�G+xq�|:���sD���&aro y��r�/:ƃ���]:꫶�$��"���V�����)M���jl��E^֕d[eRց@{� �_�o�����q*a���M�&.6�h�X� ������	|n7�!��u2��K�1�Um�Y~�+���t��d��v,��o��0L\Sr��s��|yr�}��$���7���.�x�k,I�a'�k�9z�D}tQ\ej�K_X���� ��c���8���1}'���7+��z�.��`ʨ�F�pl
�?�8]u_��t�(���.b�4/?cd��|���դ���:e{F��0oo�Զ���	Y^�ߏ�*[�{:.;�v��(��'�a ���ŐN���7mE԰|����ކ7��~�U��S�m:��\".0��|]NH�s�wY�YL���i���"���	�a�&/i�,�@^q��)a��
�=3u�����.�2��H��J�A¸�tFi������ �i��u.(B?<��o�xp4�N�0 ��0���I[^��
�0��rʺ�/w�ç��/*�,q��wL��t��W�AN]���QX�VP��E}��������D8�G� �T�� L<�{��W�����@˫�ߠ�s���{�l���{/7� �xt�GD1���K��W�{v�C��3rs�(�/��vxM�rC0s�Jf	�Cd�kJ�@n�.2(��R��PMVצt
x?$�l��O���,d'�_�	Gܔ$��S�8�畜��z�x䏜,�vy���?y�Oo?8Dy]*YlM��,�E��w�WwRJU
;)���+�}�S�h5t�b�IGG�%s�n �!�����z����%�����$�sI�� ���������kh���Yr�B�z��"�=��xL�r�@>hJ|�[�4���Y�=��2�q\�M	Sb�Wa�ZJ��?Uv��vJ.�]3'w
�s�<��nVM��Z�=ǿ��2"������/���Ľ�A��e���n�4�eɥ{]��Fo���=�3�ԣ�VK� L��+���*)���5�b�J`�^z����_1�\LN��EY���g�AG�"g�輽��rUG�&�:������,��FF���0�%'vM*Z����4�D�:�Y�]m<����bV��j@:���Ӌ�g<^��3}�^��l
�s�A��R����LNA.����ޔ}���Qf��&o�m����Jhv�I���$��ʢ�B���![P<��4����ᅪ��7A�c4�Q��O��.�5���� 2-�Yى [�g(YVN�Z�t{ܹ���A���,�xc<5�
�}�"@Ѐ��}׼����N����86W��N\k��}���T���V�'A�}�d�N��[R�����x�MEM+�#�O�n���O���y	}�]��qͅ�o�g(�9
	ԗ������"�t�Yv��2*��i�@��V��zp-y?np��O|ͧ@��b���F����Z����z��������LEѬ�M��j�MDΘ���i�*>������9*�3��b���"[�\��sNT�+( DǂxWљ��ۧ�*�_d!E9gp�pOo79 7�1�~ke�����SU/?�X��	u�M���
������f�Dpb��E�&5�� O���Dܼ{��ګ߽Ƹ2��#�U$���ZPN�M��\u��������)��LV�c��<�/�\gϴ!J���4�f����!�Ae���q\D�+ �g��&~�
I>��Ⱥl\d1��e/Y@5H_�@���!Q�Yn/*�r!s�f��#P��ar�'�L�(^q��é�.d\��@�]e&z.L���������,s7���ʅ���x��朰��"�������}$��-��%�7���y�?�G9�D@n��5#P���BK����:�w�Ҩ��=�y�g���Z4qޜ+eY�e�,�M��Ю`��rnH¯*w!�1��=q�?��U��銧�g���]�b4�nn#}y� �ڥK� ���J��58uB ��l��a�r �_��r��:a��yt��4hB�����m�M�����.�^��r@b�&r?C����L<Yz�Cf�1@>��)o�h)���M�g1
|g�W�o����s�S	E����o`��D�'�
s&��q�\����r*
�3-��[��/ft�ז� �EtX!�W+��JlD���w��,qT�#?S��_�2)�Nv��\��a�j4�ݢ��*���l);��Q�[-�BJ�~�� j�� 2�Dħ��DvH�@}�C�C%��⮋D�q�Mg��Qɺf�������+�l?!���0��R�l\�0��a�	B��T����yŖCS�!��}��V<�O쥿{�r=o���f>Im[�ޑ_48.j��U�=LW�J�щ�7�]x@B/���chy��h�|6�;��se�U]ˑ��V�^me�/m�Ԁ�>��!�LO9P[5��6���x�>�Q��H����}�� �}z�� �9�@㔥��^�1z|'�-��d�"�t9|�w�����UD�Y���+,=V�ͩaQU�~�e�U��>\yhZ7�<��p�0w�Y��I�����l���s���j�dp�j +���\���s���J:6��� ��mS��<�N7}$����bC�D�]�������-y�x��Y�C�GU���Uҟ�Z��x�]ŷj8��A}���C���o����1����/\�t�*�_ �:���hv��F�v��*-_�=��? m��������'��%.}�9Sx����;yQj���%���>+���:���3�("J�Ɲ<�ϻMi(���`��Y�Q)M�\�[�&O���z��[^�ڧ,�\=;�^L���2��P����V�Z��Xǒ1i��j&��[��.x>�!���QmŎ��^=O�<w_�˓�B��>[�Bn�~Sһܔ]0:<�:�R�(?+�0��UVJv�l��j�b<������
����}I���O���ڃ��O�[3��q��b��e�SYZK�����t4sv�K��`�b�e�ʁ_��Q�+�m��U����f�P�2˽ߓ����bLm�&��EB�>j�����jv����!�F��\:��3<?;�E�L{�1�e�p�(�Z��7��%W22���WĜ_���jp���p/i�̻P��j��}��I��u����p�"�i����iX��:v�pWrS�'��&8���6Bf`��+8��u�쥽"��)�$^�=�N�g�N�2˼�b>�QM�Gװ�ߊ�`��)�|�!9��Q�1�:�Ι�[��~r�7�����tX�9/>�9�Ic��9R�T;���^�+�-u��Tal}�]��ݛU�7>����]�~ۧ��˃[�@7����ݍ.�g=Dq�鈆�u�Q+z���am3�QMo�2� NgM��B0�&����e���o^�fN�q	�.ٿ`Ŝ�,ψ�D	<���ʒ��O�!(v3�y��̼6G���k9a�.��y�q�d����2�cH���	����O�ˌ�������ٹ��D��ч�'�y�ʴT0�T�'Z�\,�a?m��t�*ܤ��g3Ok�Nr߹�4�M�����q{^��!�-�4KU+��0�q~���zN��tEˏ�N����:�t��&�hX��b�Poʈ
P�K�)^یE}䂓C���"?T�U����O�X*�f.��C�T�+-R,	�qlbR��hk�Vni��T�!�|�	�zVUH/.��
-�I�{{v`BuG�ح���9���0T�U��e:�0��/���IK�J�R۔�U6���(��WXm�noݎ�ӳTstsl,����G���:�rSE����D;�������H�u�t����N�z�l��.K��4�gD������I��ʽZ�fIJEd��E_6�'�1+}�'1�_�Ǆ+PHp�;�'L*&i�-�=結���?���&��n�z~k�bm�8Wr��Z*��Oܐ�%eNmV��?�"sS٫_��o|U_IK�����Z���� 塱��[��[�S��Eެ��#+M&�H��ѷw��g�l�JRU�T����Hd��#9~�:r�4 �5����f�(�ȮJ�����gl:@[��]� �(�9C�uKE�v�u�^pAW#Z>����PPl9?�i�

���R C_x)�O��oE���p�?�Y�mo6Ixzݍ%��?Y���q߸���c)c?ȯo��Z��0j��ex^�:8����6�!iE���ẙO����Խ�������
e�p@ҟe(ﾤ�h�7����,�;�Px��""��#BѲ�Tz�ca�DO5��RiW�ĩ^N�|�S�5����7����S�\)dz�B�/��1�ʵڑT��KI�лk�����p�,��I|� I;@��d1_X�����+���Y�;�B���AUqW�
'��&\8������?.��D�?=�A3Fv�8`&>~��4?Ì�ʫ�˚`J~J�kOo!NJF����%�����T�u+�w���\TM��c�kLs�@!O3\X$N��1� ����"�}����/p5tA�v].*���Y�h�jIk�~��( �����$���o&U��S(�[�,��1E�dPi�
疡�,t[��� ��.���;�ĸ�cS��""let��*s�1�ah_k�F3�h�vK��(��EI����N4E�U\g��{mD�:9,t=��b��N uZ���+)�M�^�L��mʁ"{]��Rֹl�����Fd/��3����=SS۫l��yE�,�w�Q�A��h�%�8�1>����^�N"��"(�^���%,N�����V;![MkDQ>I�~���,���M���oI��(�LRD�p��`_5�c�"X�����k	R��`�8�H7ۧ���+1\������3��������+fE^�ް�OI��P'�F:�0��	�� ,��}}�/(0)F��g���?���ۃ�}�5�,�Կ�����:�lz���s��7𢝽��Ɔ��|��Ť���Gh�����pUz���O��#G D�'\���9�H�b��5!��9�7��V}cxPw3�x�;�ݐ���ձ0~��"�� Y�$;,��>�N�qc0�O#�sIJ��N�c�71M�qVv*e���;�Y5��֧�0���Uμ9��*�]�<u����>I~�E�3�hB����.��G*�������%���ܡ ��}&QE�|;b&K�Q������Y���������}�:���GnmH0�u�e�[ͦ��b�� =`-�z���v��=����E�?bL��C@������$�L�˃o�����`sO���k��=Y�f:� ��L���'�?����c�bţ��2��C���$/�� �ۦ���b'%_8�(�.g���J��Y[�G)2R9:j�%f�H+#`��[+6C;,��1Gޡ�9���9��g:_�@1T�P�5�2ևJ�Uu1mY�]	�U�0�V科o��m�Au��(� xy�0������W�;T� m-������%O��ձb���d�V�2���g����v]'l1K��ʬ,"���n1	p��?}���l%�872�œ�ӵ6��_�����8�ń��BfݹNddRvĩ��to�����N=8 D��|�ݍ�
�0��L�T&UI�V��Oۚ���(b�"k�����//�LX��/fA�L��^�$��]�%�_Z�>I�C�e:ۦi%��@ESD��tL�S@ڇ��E:v%�k#��b5.}�o�j��_3�
��_c�9G5����F/�!�����p���>x��u:����#�2Q���D-K!�Ӕ�J@���R��]d�y=Z��$-Jy����N�"���ڨɴ��re��j�܊��H���Ȥ��?	�����AP%��i%^��ع}�n���Y�����Բ�H���g�k�5 ��3o?I�0�]!P�W�} �@����R;9�i<�*>�v9imYC.�3�����2^h�n�0��C������v\���`<��,#uu%�S�� U��Vf��#πo|5abW�_V]�'3N[�ݫ���
����]b����_��OǤ�ڑ���ox����G֍"v�+8?_�N֗�x���K�_���:������I����*<�XP��E{�RV��ڝd�0#��`z��vK���S�L����;L U4��m��n =�0Иs"~P��<@IU˕=���:����	�隠S٪BR�����;��}6��Կˏ�p�����8�/�������`�3/o��/"����G��̽˲����e̕�v�W��*>Uџ��2��|}�K�g��z�4O��^�k�'��>P��7f�W�����r-�ɞ��[ =�� 'i�ǈ�$�#I�>Z�kG�L`���T��M�1�W�$����1���H��������A�����*k_�����O�0��g_9Ս�bK�XgT�|K�܈sg|"�i��2��/{o"��.[�#��C�+�a�X���R�&0_��Z�Oe�fH1�'�i}����'Y���2���[��>{:$jF�T�M�\����6�~;�4�߸IY����D)w<!�ш��i@�@q��)�v���qi�W��	�74@C�'�LZԪ��C��<�xG�c��*Dl�s~�:H���<���P�P���B#��mA���`�b$�f��т��h5���f�L(��8֫A&$&Vn���&�'�1^�t'�¸��x]�開��krRI���}�~�o�5� j!�i�w��[��N[9�*8ym2���R�뀨,��sɸ�6YBh�;�C�1�\S�+{HO}�l
�s��C
�<I>�� ��+��=�zxw[�nIW��4%��%�q�u&���?�1>1��,�����j�J�k����\H��V�1����Y
,燌&"@����r��o �~PV��#
��2�D
�Mӝ�����A�X"f1�#暱�k<N-�~mҮa��Tz�i;=�V�_��D�ܭ��LW�4~)�"K��
�"."�=�������:f���Zs�����W��D~���~���v�:E9(h���즬�+�-(�*s	q݀7�XeP��Sw����,(��_�63���Iq�Y��#��}���~nJ�x�R����Ry�}�G�$�T	T?L��ZG��ן�+��5���N�+%��4�M�F��J��y�RU�
~i��Gڭ|�~к�n|p�i��XĽy�G��l;�Y��ޔ�}U�xxd��֦tsU��	����y��5\5�� ����@���t����W�@ �yE��j����G������u�ܟ�x��e�=�^]�?��c����J,W��M' 2.�����B�/��v�'�k!�P����8���$E�
��9G�ޡ�xl{Fh���^�l��ж��L5�9g���5�h���������@���^�/�F��o����X��O�U-'�tO2�֔��M�M-{�ۧ������H9S}t0C�AD[�|������&6�\���ᴳ�i���l�#��o]	���2�r����\nr�z�iBՙy�w|��W�?M��$$��e]��d�u�:�¼��$��ј�AQL�g��9�g+����/���fQ�]�^p:���Ӥ�a�q�zE�'tX�ı)�
���1 �a]�N[�ٱ��^��*�]<��Lz���38���t����T��%�vE��|�0(C���i���9"B�\��߭�>EΞD���Ee�~J�О��~ �a�<U-ϸ&����!L�����F����7eDîӍN���!ۏx�l�s�d1���Qգ��G��q.P�O�6��w��0B�m�kt��%�����~RC�	u�r���m���|�Ў��	��J��>^F�B->���5J���&^�B��b��6�^����ٖ�E��E���&�����@�h����w$B/x�q�G��k$Ï�H-V�9dkQ*>�3�<w���	 ɗ�a&���#W��	�[$��� =1&:��lh��	�é��eoi�v.B���J@�sjԃs�i�g�kj���<��Sbg��e�l�z�����`Q=�	]!��̗)aj�뭀��'���s�29��	?Ӄ��ԾO�lQҫf��n�(T�d.�tE�6�_�Iͮ,��kJ� U����6��A�p"'�l��
w�G�3�c�x�8�>���xtڂ�=ÒM8#K�|V�2*��%?
��粵�D�L:mDSf$��FF�Pֽ$t*`����˅;���)�s�	�N���ƈ�Z�ӓ��fWT�[9c�":r�ϳ�(]�͘�V�����磚���,�Ϭ���c�sg_Wj���ot,FM!�MB�)���a�Ok���j�F��{�ֲvn]���Uq�wWe^����B�ԧ��+UƮ������H�m�GB�X�qzSrܦ/���YQ���������jg�E�q�S0���*��|���l�
�+kIW8�8�u����(��Q��OH�pY��ߓ��v_��@�MD��f��G>��k�V8�Ɏ�n-�h��Tmkإ�x݁�xBnla��A>`9;]���F2�uq��㓒��x�~����&��/Iv"�o�I�jy�o4mg�n��V�e��ҁ�ד��/�����y��%u^(������u���볇�H�� �tłUM髞���+E������A��h�M��f�PI߬ڢ�����[�[=�W+��ʗ2�����k��܆+(-�V<.>��;�ԜM;���T2z�̬�7#"v|�k6>

�b8��H؃4�gr���&���kϘ�}���Vw�Xe���E)8��z?M�����[)|;w���?�<@g���Vr�m� �kR�e��f�=�ٱ��p��
)�v���[���]��}�Gh�H����Vo��t�,�r6�Q�fȣ�.�K��n��0/��`�U��pD��徽B�TVV��K�0�	0���J9%AΩ�h6)j����W��F��,4jC�+�M-��\ۨ޶z"Q��@F�ȺT���~��hK���9�㝥a/�S��}m� �-C����D�1s�	�)٥S�{�l�k$�C :���5�ڝ����'��
�9����Q""kr ҺTE{�J����̮�u8�jt(��;Ƈ�EY
л���\)Zq�',,����|����Q�5y"�op�5k�꒧�ȹ��<٠䐲��i`f��I�hS���}����A�c��Lǩ ����֩K�Nl��\�*��m���V��L=LV�=|ٷ���@[Nm�pM�2Q�w�bW՚�<!j��<� ��-�KNw�pl�����b�`�)���NO��q�U_�>(����d̀!ޚ{�rʥq@jZiG}x����������dK� �k��g�Y.��2�cGb�����]v�;��_#}���.�>;��c,�S4���vG=i��S�n����f��a=������<�t��rN�FWʄ��W���}���W�o�h�أ ����(�{�h=�:�h�����ϙ0mX��}��u^��BDī,	:�GG�5U�|sx�M1��9�������Y�|Ο����D�,vD �GT� �)��P��W���7:��ƑY�S��l��tV����q>T����t�M7́��t�9sK��o_�+*kqT?�9�~�j媮ʂ��y�pA�Ê�J��kE)ȱ[�h�,uD���ba�<?�$��g������T̛�)]T���?�gإ!�:"\�,���0�J��9��'���>�>k�k�?±p��{i���:�b��������Y�����l?<��3�2=�� ��׀t��ѥ@ ��ѥ���a|;ϥ��e��2��2;��{���k����ki2���@���yqV�4W&�Dk�վF��(b�Y�~(�|�Ry%H�ޥ�;�~����2� 2��yf��J�I�N2�h��A��=���TI~P	����-�T��t�>̊��4�Rc��g�4�[�[����0�@�����)�f��}*7h�uWa��.ꊏ�6`|7nR	��i����t:>!�Oh��Y�lx�uQiB�׊�;�C�n![w��jc~���I�M �h�b�u���|�S��8�L��z��Tdv�|�W�y�vMV��Z�)!�*���V�J����e.>ͽ�8Iz�^��g�/!Å$���o8��Y�BB� ~��e��_�o��3Ť��l:�V�圻��턑S[�X���_G������h���uAI�qmok&��H�\�$���T��%|_��̌��x�G���+Z&]�׋�������y�9m{���bܛ2>K6��ʧ!]�y@a���*��4��D_�N��E�) =z��,OQJ�� �}j��(e0��N��u6)�M9�����y��[�8�/8�掲�_��* �[����]��F����OY�
�u2��I��
<��,�&]�P6� ;��'���F����ˎP:Q�L|���`,�V]�0s[�DW�5X�d�r�,���y��.��W?¿���=\�H��5��=��F,'�"�%�C���J%.���
�K�⫈0F�Q�TKK���t5ty�Շ��<6���e݂�`���h �q	�+��o���G�^򜂍�=ݞ{���H˜�ȔĤ���������:�~:Ynh6�k+{D��ւW�[�B`�^L^ѓ.
Pz:���g�{��F=�#�§T�"gU�ٮ��v��@hI_�+�YqԳ��g���W�%�Ծɻ��r�e#�Q'5v)5cqj~���F2�o1(#Ta@P�ѧ;��⯯�E5T�P���8,���������-Z�8jn�6��y��su\�OK���E��ZYnϼ|���)�_Cs�& ��Zل��������u>DW��1JeT�)x�|�߆���x m4��:�Ae���nyO��0��� %Z�U�;�ͺmُ�f|��?�����[�?�p&|��P�V=8'�:Z�6��z�_� ��Z�D��s����������'B>� V|�Ӟ�b3�.��װˏ�LfW13!�px�M��EǱ?N�
1�������{Ҫ����>� S�q~Zd-"3h]�9���ƈ��J�-��\m�`�)�M�B�5��S1F�Y���NI���+�w�>t�����>|v���?RS���N�|9���6�����~Ǽuғd�y�[��c{{6�O�7�On�n2^x�f��6�T�V��y�A���(��礙���D��]���0���f�J������r��UI����E@x��dn4�&�`9�K�$M�-��O�Ow�eg;p�Z��� `���7\��hx���U���px`�z�!
��Z��4͠YW��Q�P���`�5/.�}�������q��i�§'y�s�(�� �)��F[�\��ē�g������-�=Y�7z�+-V����flU�����\|��{3-.��w.�u���B��i��C&�V&�����%��͗���G/|��+R/��#[آg1ޙ//�OM��ٹ��(��#���N/ڼ�KV����|�D��䓭�5��
(���	-��zm�
�)������,59pUη��F��� �N�N���}�Q/S�*�0}�)o?$�sX�0-mRם�ޠ�S�;2�^߫�͵pW%��͊8#��0������Mǈ�e�,r���dH�9���u�,�-�y��+bN�8�+Tl5R�C�Q��v8�fP�?{�WSG{���q��#�y$0^�?*�UmΉ�FM�q�?�l��}T ���]��a!��Z@������Cü��<X�������7�^���,�7�`��y�����\N���{z�5��r��i7�Cygō`������/Q�`y���7r/z7��b��q��;n)�d,�1��1����@f���6��$g�.��@�h��0F��`��]D��ʍx�Cae�7���H�O���{������N+��%?5���y*w�l�n�6���-*4�1Ig�w2]��?]?;�3��9�:8�%^.��pxv5��H���
��i�E�;�����X�.��$�>��|x�=\w)��Ap*i7O��≣D��D�jI�/��0%����w_��E�3�
*D��Ms���ˎ�m���2��'�TK�=��]��B��?`�ȗq���	���W�n�|Dk���
��"xG[��"s9  a]nQ�e5���ӳ��Nn��9;����F�+��gΙ� ��ő��cqʁ~��/���ǝ�2��O�b~�$�� ��������V,��Β��V\W�49] ��ZY�M�ͪ�P&�����3���oNʶk�I'y�h3����{���TU�l	^w���X޿�s�.�-��+(P�'a@L�b���1��(Ւ������A����H�O��6�O`	FO\�Ȯ�����>Ҧ���M����q(v�C�?��T���(��E�Y�j)(�j�:�����M��T˴-�t~�g6�JJ��}$�u�X%<�N�j2{�,�~�VgXTn؊����r	�1mR0Un����M'N:k��%P0rM#�B,���3�\e��죒��o���}�����7��*ֽ�W�����^߉�n���z��_�Ͱ��N�Ӓw���D.��J<G�_>>�Z��顾\n��Іr�x �<=��,@NK���M(C�w:]�Y�ϴ��)�"��Fʦ�|`��T��NCTyV��Ğ�?ۜ��#kZ��	`�""�ߞN�ͤ�AފX�),���ù5K�H�VƠ�:��k�Ell/�T�+�-�.d<���ͥ��Cd�7*l�_H��l�ڃDQ�vH�	z�_��� A�Kr���qV�`C�t�'>�m�����j�%�=h�y<���#<J-z�_��g���q�J�٠�<�)<w!�?�Kw+0��1yT:�I�r&��_7L�
H������I��c�ٍ�1��]�����.�Vx|^��RِG0%�R���""�C
�l;�L~�s�����ֈ�k`ra ލ,觝gG�R�8���|��E���̾G:�m����"/�;x���^�#Y������5;c�������|7��Lؐ�.����gk�F�
���g�:��>F^}�gQf�v�]��k��8�/����߂�����Z��.H����Eļ�|D,[��-�|�
S-P��t=�D�/���_.��`���7	Aw�)웨��ʵ�2�ԯL�'�.�X����_;C�=a�z(�P�
3Ƶ����}��Z��!�m&�H�n/R����TA�>�q�\5��z)���n ��F"���>`��{���)������.���&K���3����l*��d��O�p���4��Pߵ��N��f�Ԉ���f��������^�Uة�"��_ІH�T2:���;�7�EEh3b��@������Ġ��7x�~mR������'�ȷ88��AK$�o6�\iM@n�ݓU���ʭ����b��ĩ���`7����b� tJΚ�`�m�|'$��F��5�4�E�,��biw%��k��O��mz,�EN�j��1a�Ƶ�O�_t峃�%Rs�/ˣ�@ѳ14�Q�loh�٘r��Z8��{���-�\\��-#���ԐI���bX�s5؋q�g�e�"܀�~m��T1q���f�y)P����5X�d���I�]��a3�8�c��[��.��T���uS���}X��+��5@�F{.�0dD�.�go� ���%�2�W��^
6m>9X�SR�r*�E� �0������T�QK����]=��ޮ�)����p����Э&�� �����͔�x���yTQ����q�yT�q��vcI�)5�-_���/�h48´��l�C������$AX@[�}Rʐ*`C�π�u9u��[����Σ�H�cw�X@�r�;4ɟ���Eg����-\������!HZ��XCpə�ɚ��E{���ݫ�3�d|�ֽ��~/������X=��7�{�wJ]�gC�Y�ݴ]a����e�4��ފe�7QDn����߫f�w_lK=$+-�.�'�'ؒ�Ks������
ay�L=�1)ٳ�S襪���y�7y������3�"g���V�䆙�P.���YE��8=�\r@2�W�R�?l��N�P[IۑB$h�s���Xi [C�<�ڳ /~�,� �d�"�b�8�2""U���k��'���u�'5�毜�	֑𿅈��o����1���)=�x0�6�b^�{�����,ғJ�n�W�Y�X��>�p�U���|��3{:$bz��{ჴ�x����e�smZ i���t1���4�ʵ�*���i���<���2mI�߿���˿U۩���1m\��;!�.sN������k�g�� @�}�P�������?Y�|�r��u���_�of�&%�F�5|�����l�3D+�o��0���L�ǟY�1MZ8��������(�`}a=s��q��θ�� �>��ģ��bWé�ŉF"�>��|��M���K�җ��92��
f��#Y��Q�?�L�"�6p�D4�8V��y��2�Jn}x��t&�f��7;p�$,I+�x��IK�e,{)�:�z�6\@��OGs��K�2i���}�:M��G�]���u��Nb����;��! ���q� ���u���'���#d��]C���'|���y.dv�Rc03M6<�j����J�'���l�]J�o�a�!g^.я٬��\P�jz���=�Cn�^CԾ����3����O�V$F���&�F��фѴ�(�x'�����H���jHd��k�ҕ}�TO�t�L6�A
F��61S��2{�Ն��R,Wk���DM?%�#�"e
�X\1Y\�Xc��ټ�|���e�m�����}}����H���Z�ӑւ _Ѫb��N���v��C��_����
���S4ݠ��Ft�'��nG�����:e�;]I��K�ce��(e��Q�7������l~���#��ʨ8���>���qS�����G�ab)�1X�^G/&`pJy�9�Nr�zߡ�4 ?Մ^r'�w�L�D0����8U�M��g?u���U�#�c�cJMU����[&�9ON�*+.  .'���!Dĝ��f���&&�K�!��O��F�9HoQ����{^M��������;/%!�)�t���^�������n���DZ@�A��x�������p��=g�ךkνϙW�+w�t�i���گ_�A:�_���ˊ꼿K����3I�W|U�8�x��8}�#��eB46(����
}�k���U
��ţ�5@O�/M̝c@���Q��f�ܐزf�}y���*�.����gy��׿M�h�d�%�-���W⨛2D���P�?�J����v�.G'{ps�w�r�T.�x��,�2%T�w��(�yP̐�U3�c7ޚ�Z0WH<�xA~Ƃ���y� �A�l'D����'�3�dd��?ѼyGM%C{H�1��TN딷�]��2�*f�*8J�5$�fS5e�:��a}g��}���Ҍ*{􆉍��h���wMA����k�WM��~����.	�����uyH�L�0���'���p�~���q�2��%�.�*���GUT�a)	�$�>��#\�j���S1%Z��3q�P@V��DH����~�����|��+xo�����/��H�kY��\�Qugqx8)�^Fg�ٱ��N�%T�6Z<0����!�O�pb ��w�x�*�f�Z�9&��+k�="󓭬�duy�b�7�9�!��Z�* �*F���[|���<ωy����י��{?f��'���o��'w�(t|hJ�{��S��H�܇HW�O�E��:8I�b�@��!��t x�C�%�%��X)�W���*z��U#�|-�sV���h�yo+�'�����?V*���d��������m{5J���GA���r�Fa�{,U�S���6�t)�(�i��&h$���@��!$�i�a���)�샓�I���'U

t�<\e	�m�^�	�}�#m�u|i�ѭa�qM ��虻�q�Vu���a��B~�
{�fш�2�����ԣ{�Z���p5G��n(��/]�#����ۗ�n��I�[�=֣���L�^{���9Pڰg�k�aOHu���
O�E��X�C����U��Z��s�;�9�a�<H)c��mY��3|
e�.�I�`W4�tx�b�F���s�8W=;�c��r���&�^�}x�sa"]�`�aR�{���x��y��_������1�H�Y{]��侓/�����OF~9�i^�^��kLLR�7ɴu�n�?�;�B��T���r�i	�#�G�&�+ :�m)\�2��	H��5��C�TB+r|�|��蕆�(TB��|<���Ս���`���!c �ߛ�V��֬���5/61c�e������N.nPM?��N����X�+�DH�8�	�$�����-���l�}�8Hs�\��f�7}:ǠW�������41~	�"��}}�AB�3��`�X��@�:Ф�m7����,B���HK)ưê���$�Z �"�@x;��jۆ�|C����)B�zKa/���������s>�ڼ��_pS>D��Y��������%cnҾ.˔����!�2��-^�T��G��ї�A�H���n}����V�	��RMp�J��܍�d5�?�������?�����HN�-�[6���R�]wç����#8������]3�d��^?V]��|`QM`��RE)� ����l�[Ѻ��6<��&J�2���P���/Yc���sO�Ψ�P�	LF��I@Rq�\���#���H�0����c��Y[i�e�F����=�8� ����ٸ�m�Q�&�(�.ӈ�],�Z?����r��`�B� �BI+-�ZS{����>v�3���&h\��J��M ��0-ځG���Y7�u�ö:"l#��BTe�0��ոQ��@�?����z~QL	e(��v6t;ƫM��"0����T�Zƨ��5��;���`�kD������v	�;��x$�؋�Q��NeO;�n��QO����1���
o�64� ���!��o���td
�B����,�vn5�ވ';�`�(�D)�h-�+h�l�$]x�$@Z��!I��F�3_�iѾ3 p=�G%꽷� �A7X�k�9\x����=���[D�Fv�����/�c/�D���p�"����lj_�r>�,��]���#���UN�8���:9!��,�~DO�ㄽ���8;����
y}�����T�3�X/�b����[��/��b�]'�^��{�P�I�~����g#����դ�L�[χ ��[���_��b�ݒ�A
�⑭_�O���r聾�����&��fk�K��t\�����+�����6E��P�0�`�b���i�����-,���)���ϔ�o�ߡ�W�f�8
<yu����m��+;.����fO���N����*2D�'`����ޡpVz��Q�Z�U�w���y��mسӖ �5��[��C>�����1�H�۠�/R�A<j@@M�����d�F�C͇��i �Ko�C��䓤�{ߺT�W(>��g�T�,r���?�՘��SoH�imC�`i�
���P��m'��n���򪸸s�Y�MW���!q<�a�w>��m|�t���@kp���/b�d��xYOŇ;��_��$[
{���zcWwÇ ]Q� ���g�\�Ez�ls寵�s ��\v�a{/�Kr�/wL(�r�f4���+=ع���3��O�N2�f�����,��g�A��.b����w/�5�_6pWD{��--�1�em���q?�ւљ:j@� �m����!�8��y:oa��+��|�(�О�C���K�|�ZdS�Q����>dU��ʻ���0��T��L�X�ț����f?yB�-5?E�F�$�nWI �S�6�s�}Z"oH��3ym�hi��=`�v�Hlj9�K�K��1�W��k�y��*D^}%�2�
��� ���O�H�i�������p�=r+G��B�V�a&�HF�����>ȸ��9��){!=*^y����[��
Gt9��|�����n��w�K�9*��;�4Qљ��
 y���&<@f��0Hz�MtF���3��D��p�?�X�Wq��þ�F����g����E�Y2��GҘĆ��嗅3���~$����������ޫ-4nX݈L�P��R��(|%�2�Bs�R8���p��mq�R���7X������B� ���b���7�-�/#"�$��.cW%{��	$��lf�0���y��h��P�|c��C���h��I�{�3�y�vV�~�&��ݻ��CȔ"/�\��� �m�|Bc���$�.��z����?�Fw�
�ۯp�4~:�1�@�c^m��5���(7��2�_G����jH
T˫e��g����?1����{T���/S�B:�8ѻ��W�V����t��Xe��m�����̴��^8���4*4���v�E�[�R6�c����~,�k�Q�ۗl\� ��y��pX��T��]��`���.>Q�H�`�e����6)X�uQ�o��0 �fc�ƭ��J �|��pk^Ϛ�`6?i�i00#S���00��pg�u3�~�~fv�����V�I��b�}4Ѕ�p}+��2�o�d�޸�s������W�q PSc+�#Y�iܻz��w�O�V��d�d"�2�G��L��j)>/��6X��hϝ�(�R{�|�������#%�Of8=c#���}X�ضx�a�<�� �yY{	z����~�k�� ���|�m��[����r��G0eb�ޤ�+���H��Bd3� >��9�X:�L�Ӛ�R��x�Xd�y��c�N�U.%*C$!����?��W�ဎ���$�c7 Z��Uw�Q4��р��q�qo=:Vq(/�,h�9)�X�S>�B��J�[C_��fH�h3+���-h�i��ړ���C��m:��Ō�����M+�6b��49�L3����sF/6I�PǸ�e� �-��G�r���&9��*)�>;��	@���[��򋈮�}�; 5�m9���ä1�&��:��a���V��8�;|U�h���78�ގ�X�B�����=T����p���~W�jߩ�:x�}��������JɃv��%�97�^e���������70ۣ��J���n@���1���qD�&���'�#��r��S����ti�A`�a5@j�%\���*��Z�D�I�7W�(b���$d8�e�L�Aݨ*LK�0^Ln�K�nL��-W�����a"�Đ����/G�ʬ����"εJ��ݳS^� ġ��H�)�(Q�Փള���Ȅ�"�����ٶ��5�B�e�M�3��s��q�7�`਌��e����J�MA*~�B�F���=�f��k�<�ܵ��?��n�gM��_�.e��$)u������NF��.Gt蹰1U��.Ӄ��o.m0
�dt�#	�4I���B@�6]�q��*��+Ԩ�x�&Vf���;�����(c�=����ܦ ]�F�����x�ѴM�0�4�S�>[�U4�[ nm��v�!F��X�3y��-ǔϑu�z�h��J�ϼ�� �)I	%m#C�I~�z�C"�Ҏ�����1_��'��N�T>������4:cI�ڡ�Z�m��Uͥdl��Y��X$O~��^/�-�.����{��Ǡ�n�����{wFL@Z_��c� Qb  [2Wo}�呶���L���W��-�!� �V"�uR�2�����g><��	p�)�*G�'�ad<��o�iK�� �Ľ��K�_{�2eLi�TV��?�y�����$�D�<�.����Vf�����H#�o�9Y���\��L��״�]
Ue�^�":-g����,z�kuq����6|�;N�:3��")�/��C�4�� �Jfڮ�;i�����oy^"���&�y�� �'�Q��+vI#u��_��S��k��ʮ�d?zS7��+
�Yj+ĳ�\�� �`�l���y�2����,� �	���h����vƞrB�0k���������^�
���I� y�C�(����J}ػ�J��8?\ �n÷*S�i�P!�S_��� ��vj�O��q��$i� ��=��JM�z�	�.�H5��>���I���R�U-Wh��[%�AP�Uw]=����"�߉�P����Ͼ��É�}�����w���*<�-pOJm���LW��
��u�v�T!QkE�rLԀ'�����9���ѵ�A�C��0�Cง{����Nn!,�2�c��I�n���R}����Q���\��4����ѧ���m�Ǖ�9�h��z^g��w�=��J�E�;�${)�!�Z�u����4fbB}6g�z�N���g��6��q"�t��@1���biB�a/~vg:�L�Dk�L����r�4	�i9�R�8�5������<�6úC���+���d�C�=Q�9�����s}���}-�Sk��s<j��`��Z��TY$T3s���`�t�+eנ���*�>d*�r
��8���G߄/�Q�up?���ely�ŋŧ��$q�xȀ�8�&��l>sI/��v��|��@��G�m�!D��b��a����a���jJ�N���φ�K췭��|�=�YQ����[䷓/�9uk�Ϟ-�=Cz�����?+�����]�w�XV5��o���r�2���jR�oF,�L�I��X=n����͢���s��`����n2�4�qE�(1xAm�!��2�{N��eoF�	K`�2����pF���ّ��������>�lDH=�f��p+�X��'�W�(F٪G���{L���e\����5�v�P�g��k�:��~[�9y���w�V�����3�����R*�&�br$~���U��x����,���'��떨Ҵ@���DH�h��#~�ye��T��W���^�xeĩ��W'�$䱡R��3H�LY`�hI��}v�"}���5��;N�1ƞ=������d�H�9�R�F]�!��x�5ܯx� ߎ[f� 14��'��'����]��Z��K�%,����$�ڔĮ'�xNmGE{n���:f��Ag')=�L-�U`c �{3�V�;]I�K�ag��>�a6��b:�Cb�x#rC�x�I�hnIV�Ͷ�B¬Ҷ�lz��z��%x
�_&V��!嵎pF�E��5
�$$1]q������!}}��ħ��S�S-��v��j��]ܴ�?^��RǴ�+��5�h��i3H@���	�,~ML���@+���xhRWz��C�)a�f�j�zu>"[Ii��!�6~�}#\!�*�g����p��v����1��6�� hn^{%�S��У��R���
��l��W����"Ǻgy����^�)x����nf���s;ː9Tw�A0������޶��EY&_o�O�PӁeX�loϤ��׾k����*!6Kf�[!�]��fQց<;уdU�fD��E7'7+�����ܤr����ͣ�zCU�))x�fKиue��$�jC�)!$_���ȇ��%�S�%t�}�#:u4v�M�d)���>&
�ތ%ݩ��[r5����Aژ��;�(!� V5|.��$(�������h ���_�s�ǈ|Φ	e4�����?�Ed_�6֐|�j����Z���c�ZV�����ot=��q�ב��P/�DO&ח��UBa���镐�Ѡ;��:a!˭�:�6+䥏���Џ�ļg�h�A�>������.*�6n.F}sb�}�E���L0s]OU+3+}H�2n?��;�Z�M~���4� ����,�}%ߙ�������5�Y�ѐ�B�c=R����<R��;k�lف���!��#�#�Z�~�C:���ӂ�܊R<D���YqBn#���o0b-]���'g�ӡDF�ML,/}�f�w(�}�h�fg�Z�����<���T�{���6����M�� ��U8�|ȷZ��È��9͓~�֭��i{*���HiɑT:��6��k�[�������X��<��b_�u�:Zυ��v��:��(�&�Q�$V>���Zf�gav̟kk�f�!?\U��E�)�\�)<C��2���U^X*g�X�͋���Z�5Ri�x��\RR�?
zs�s͆d^տ=��q��w:��E�S����A|r�YJ�xU���,�SJ<���ղDe��t������*�$D�i ���:2F�E�L����IX@�Cu`Q.{��
yѷ�ݓ�}�;��%ܡPhn��^����Bfs��>ȳ�r	B���4	̴'j:h����XSq��������Bf�Ӵ��5��������Ġ��sTD�[��O�o�z�OJb�;��e&*�Ӛi5���L��ב�z)�n�,F�):Ac����8_�i��������v�/��1�jD��k�W����P%!�$�ҋ�]j���M��]��Q��7�:KI��o��T����A�o�kl��3|%��Ǜ��K���,(�n���NGvub6d]ʭ���&ҽ'.�]N��� �ly�X鵮K��v㊰�.^�b}!Ǎ�L���=]�0��ZA����ʶ�fC[�E�m�}���-߿�����l��T�ӛXî$o�/��sm�pc�TyJ��(pR�D��H�,�F�r��������(�Qb�s3�XÈ�����J7��X��$�-%FQq4o/�~8+P����R<�\%����p4�N��`�b�T2�TR�.2{��tFodh�..�c�Q�?��<�NX;z�9��B�YV�JN��$��c��c �u�7h�xQ]^\<��¨8�T�����Hu��DG�o�nDT|��nYߨ�#�k#"r�8�XΗ�b�	A���ڂG��W���TtL��jǪk������e)2l�d�͢���VH�����[�c�\�99�dв�z��62A3�E�
Z�^��ă�5��I��I	��D�J���O�����V�j�s��J�NnudT�PS��8��aE��̜2h�3B�m��n���i��TK��ᦑ2�E���e�H\��CУz��Iu�~}ʺ�^��O�Y��{'��a�L<�<�%ͷ�������gM�U g=vi�d�'��7&�֋�Ȧ�|,�4��O�3=�el�M+ʼWZE"��]u,���t��o�%�׽:�,y�(�v9 �qHēN�P��(�eŽ��Y�a�.�Rr7��'�v�uZ_q}�����ઔh2�<E����׏���i������@�Ġ����!n��1j͐�q��B�J���O����5�w�z�ؗu��4/��"����߲�	�$�fױo�xg5�-��2��6���<����F��1=�6c-9��Ϟy�G��U���Jd&Y5d��	FBXa+:�S~o��q �yT�Ή벎B���x~V|`�V!����}��wh��������E2�Oe�؀���������)*"l��n�:�_D$N��ԭ\��5�(���+���$Dt�q��F�.i�T�H�����C�h�5���eF������!/Ny�f?�O���Z�d-v�D�|R�-�ui����$X��?��9��6�£o��q�f��k�����s��_�������Q��~y�rƦ���_ekn�S(�};��� �K�SJd��m�6qp�X���DC�2����Ȟ޾�B�)� �}�S����<���n��:D��@A��#��uz�N�{3��Y�"zx{~�b x� o5���a͐Ђ��6�+��5�b=|���r��0r)�h!�B;���lC�r�7���\�d�a�4.���t��t�3?r�7�g��P��I���עaʶQ�앖��(Y���qx
!�����
���� D��0�°اYZ��1�`=���4!�c�H�Ur�V��n�tu`�g��'��|�uQ�|��%������l��Iu���kn���1��~��L|k�� HK�Fv�ԗ_N-��GYR�J�_TN�Y3`AU[=�-�@��ٻ�?�P�B`*�������!�!�C#ا,��=G.�*+�5$c�^����
�T5a�~�I�����(�����8�Q#��#�Pqwǧ)Z����o���M��{����aư��Wy�s助��tQb>[���1�a1袓��0�᎒��q˛@^�~�1{�2���a��8���n�R�K�	�n� �?�D	d`�����������p�Y�g W��
p�u�nm^&�{�� ��|#��@�T��!W�=[��Yxۼo�E�6J�i��j��oy��a�֡��`T�-襝�G{���H	�9���%D\�g-)�H�����D5`�+���m#ݯ¨�����
�?�����Ũ5Vf��2��[��R>�`bu�S(��g_��O-��~�nz������~E�I����̇�o)_襱�9��~Tvz��zx:�y<�]�����=��t���Ӧ���H~���r(�P1q����ױh3-����?&�/Ɋ�H��s���,���Eb ����OCP�f��p��m2r��#De�̰��&M��2za�	���W�����U�۝Z�8U���Y`����YKn�C�g5E4�_5�8�$��"' ]؎��F�:"�+�N�EE�Q�~m���.;�N�`�`���\����Qx�*6 �|T��=��m�'}?#����X�>I�Xj��,��z�~ha�Sx?XEO��3�����1����
e�``-Dx��U6����	���1b�l�p�q�)2A�&]�F�ڂ̖��Z���8(�;nc��)��d���sd��}�׽j̶����`�p���-Km�Gǟ��%��@]��X��E����5���&

�櫛�l�Xi���������P������"�b��@���N���kG`P/w+4�f��eJ1�K���� M��@���(�2B��Ys-�3L������������ �ٹ⇵{���l�l����:��r�J�� �%9������TCL��0�a�-@%�z�Tn �B	�3��ى����_�=�)�����g?t�K��x�m��.m�V	qc~��X5]����\=A��������ݕW¸���f^����W���]g��@�����{':�<���	ߪׁ��� Ă�h�, ����إ_�e�}܌����U;��U�"��]*���D�NJ�m���Z�'(��ڝ����"X0VM1�b�B�a)�㹄���"�)����6J4��XS��vdt�(W �UH>�5�0S��
��Bhl�Tv���@^��8�vנV�9����������k�	�n���}���J#��E��6�&JX("��Ur3)f��"�d�X������q0�PXXq.eI���٭��EK�iT�h�Rz�a��zB؈�q�������C�;_��O��τR���+��6��]��2�gvA�,�q��AN
??�� �
�L�߈�����}��>�������9��dd��d4	�噱�Fl�w$ˀ�߲iT�)�7Z�hr`�^	����oDG~R�Kv�%C�@D������D�ų���D����t��h����%J�a^x��ZwȮ��?�>�̒���sf��\�#����L�D9��_�����B�p>3ƓVc'�!�Oh̨����gH������E�f�C���G`n��F�6��o\}�$�c\-��5�n(��e.������cvuB;] ����Deq�m\�����o�rɱ<x$���@v��=r�\�����>bPb"s~���5�F��Ƃ��?-j�"�	-�"?��ڇ^������f�_1f7��t�t�����`sl���0;���5�ĳӷZ��}�RT���g��I�E����aJ���1�7!,������vQ�⧘726��
�Ϭй��BԿš���z��Ź����&�­#�\��tK^��?���z���t�N�b�+.��I�h_��o���0��N��"4+Z�3�Tz���G/��@�"�lJ�(Q)��'>���3� ���i��7����7�ˡ�$Y�g����^>3<c��w�y�p|�bj�M |��TKO�Z�w>m@�z��k�8��J��Ba���|���V3��X����$c��lǜ#�#�5�z���I)���v<��?�`�q�����@�7 M�2�S��Zz���T^I;���9 -U̡N��y@���V�#���}�R}50��3� :�D^	���B5�j6.L�T�<��,f�� 9�7�0�U�&��!E�
2�V)~�VpFN.'Z^x��"_��\�g�3
��=���­�{����7l�|<u����x�/�ʌ`G ZI��X�_�<�c��Ѓ�EiN��Y����<p���+#u�9�V�0� |V.�5s�ę�L�w���RΑ���e��r	U��CU��I*���^A܁��F)��1�G�ُc&8}tԟc��$� �� ��1b��Y^����w�@��ƺ���e�� �h�S^� t�Vd��&[����le�(R�H�I?#=υl<Y��
��w�:�D����^nT�n#"���:��:�i~�Ȫ�Ppq4E>��ˣTz�:WF;�l���.�ڻ�H	=�0�ޟ c�-��m���9���"�FeV�y������1����_�VtG��̣����M>K�J�[����= ^��~��k	���(&�"��N���6*q��������JF9���W�uA就��g�L����Z��[�f>�����X�Q��Id��<�&�]�Uz��2�h�=�� ���3d�dTܤ���j�"Z�ͬȜ<
5��tb�0rT(Ɛ\	����FY�lm��x5K^u�� /Qܪ��F�|]�I	'��յ�RC�F��wv��*K�6B�1f(~;ι��E4���	�j'v�M �8)��w��|/`�K�%�L�a��QHS8o�͘j�%��y��y��̂�~ �I2rŨ�K�\�0���7�b�&��Ǉ=��N5q�-k_@y��aH�_��8>C�C�7L�"� ��%ڀ;|J��(�F�W<��P�8���g����CC���4�rؓe�c[<q8��8z�]� l�=�������D����YX�t�8��=M��N���6k�\׈$�.�α\�o�%0aN�ߐ���-^��p������/���5 ����\�~�J%#��E!��5��%L;����
����-,���  К��y��Z����Q:���ʸ+��Ȁ0�3mH��EP�&Q=�p
���dB�pX����,�s���\
�ycN�8YՄ��[��Z�z��䃾y(/�L2�}�O����J�P�d̃�C�ja��GW�|��FD�ն���ɐ��h��Ƃ�	�Ȣ�e�� ��D�������,�H����a���~��z��V��}������z)�=~��Nj����Y:���x.��m�q�|�O��؍?���Ђ*��[�<����!mP������w��v�A�x7V�����$����Z�exm['��Y�A��n���1�Z�D�._Z�tJ|�1�K\���_�}\�a]Y�0��.k:���(��L��GcEN�J�(ϾYยKE�!m�����V<��ׂ>OQ�Si���������&;	�oJ�����J����n��	'g�Er��+z�G}�;�(�W$xx�is7_��8���CJQ[R�'��O��K~-!a}{��L�a�%�͜b��G�	B�a���h����;�\?ˍ�Q/��xc��`I������V���@�nwb��vtU$����DGBm��/U�����M5ղ�o������%h�~��ͩU ��w7��O?��g	y��
b��ʋ� �� ��v�K����E<�̦�Bm��A��9�B-@+vJ�"�Íp9�N�Yn�u��;�x|!������P;NxW�w5'F�3�����7z?�N�F�̐o+�-#F�6L��CuC%龕U�+�)A��{��e�w1)�Ps�j��U�-vSB���Z�w��s��@afk`}F�i�+�i��!ˏg����M$S��RYM �5-m���:oֶ����W�������3���e-2cdԣ��Ϋ�tβ/Y�-�s�ǿ�s���QN�Ħ�=Sr���H}@���}_s���
b,���a%;~��:�Z��c	�|��j�m��PT�؈��'�5�x�, ��UUҢ���!>�f������[ �Pw n�J���է��\-,k�F�����8�[�A����<���v!�oaPuMCR�]��~ɎR����7��!|�拱T9չ���/�e��[9��J���U��.wm�֢�bj<��^p?��X1\Hy0w�"�sv�x��
�	�{�/_-���E�����=���s����������0�9���t���D����˵<��XA�&*%U�G1\2����1~��.���K�B��d���!]� =C�t���%O��y��V����*�q�S �6�h"�)��_����ld؀9t�*B�I�ه|�?I�w+���*�^1]�!�ͬ��N�.g4ׅ�i��\���3����d��J�D�5�7zP�Z�+d�%���+��i0�}�V��7�oz����P�(�dLG(x�l%$V���k��]��k�t�#!�� 7�y@?P��#	v��7\� �� �
���N7b�C[m��ڧ;�+�,�;�}���j�m����\��lϸ��{O����Q�@��g�'Ip:߄O��k�}� <�Uf@i	v�l/��t&Yˈ��B�]��n��b`�X$m�a��o*�-� �k�z�U�Pۙ�P��믻��s`M㑮۲/�q���д<�8���U�¢x��6����{�P���'�kc7�Q�տ�( ��_%���N��;��r����T%�X]y�و8�=P�rD��������� U9��Eba�&َ {�2��E��<A{�����p��'o�Mj��^5��L�B,�����ﲆ���WP8��D+鏮.���=�t��v��O1��>�z�Μ�|����+�~���B���*�"�=x�wΉb��%**�Vq]60PP/�F�(U(��I������Q��0���0G����^�9�7�'��G�k��Uyx:ldA��~P�Zw�
b���.���릥����Sǟ��UG�ZC�!�[S���h6"��������1�n:�����ߙ<��8j�u�s�`�������g��N�+A�0r�ru��ԙP���5毱��	���*��}b�XB������r����⵫���,��Yx��`6�`S�]�6�~[��E;��=Tr��!�v���-���Q��U1`p�@�o���CL�h��3<0��V '���<�,�Yn�U��ڲp&D�h�!�	t� L)��s���D����O�y%��H4`Qii�f���]͒� qc��y��{ԍg	 ׵�}� ����~��Zz�}e_�{D܅7A\��G'.��|��S� y�O��fc�O�窣���
�����*uXU��12���JU��<��'�{*�=�9�\/�I��+���F/�B`��'�r��(<e�Jc���.N&�w���P6���S����ʀgA�$�����O�����Qǃ���� �rV��@c�Pum��@0ё.��5�P����XOƒ�9����¶\�y���JL��6?�6Y�2��xU����q@U�
�<G��e����}��!�3�xܐ���.�^�Dgg[I(����"���tj5�s�QY�y�����NXx��!�:�g,���%˽�5%�!���->�s��D�U���x�Y 'l��o=+U����n���<�}�i���v��4�ߜ���U �����X���U4�n���F��7ћ`E��x�$�?>����D�_/r��1{�B͍��%���X
Y���Ŀ�H���-�"،�N�ɿY`����i=8>��{��%��&9nod6�g	���(�%y�?���߾�G��ױ�1�8K�'F��q����";ӺYA��􀵠�T���f��Ә�a���X��T�e��
����Г`�ֱ�qf�P���^�����KЩ+^����7���h�m�䂵�(Z��"�}bP�w��!��x����ςP���i��W��	�����#�;&b���cj0��q��nX\Y_#��%N�2���EY���$n"�6qF�1���=�4���u��$QTf�(�_( O�8�KGj�+!�OQ=�/(�x�9d� ��q�k1�e�����e��PĽ�YyI�+w@N��8A�:�:F6{sl��!��aZ�g��[�5^t��|���DU�AV�@o��cJd\�}�Ϥ�� +%"}�#q�7�un�, CD �d���d���@O���(+��$g�0#��J\�ղ�]5'�S�c���\G[.��f��dD<��1v�ߐ�m%`П�W����؁�����߂�������M/�A("����V�)�)@r�k��&�C|���bCa;^�X��NF��<��1��/0�y�Zs���C��7����2����}���or)82��~����p�n��$�����)8c_2겦��+�����Qks��r�
�e�bz�h$��������#�6�6�k�X9m�3���m^�_���}�{�	^,?_��"󡒴�&�������3��vv��N"#��D��=eƍK�8��y�c�-���
I ;���z�O��}�~�87z
_� )̏��D+:�D�5\C0�\���~:jc��t����,jR��[�����g������o���P�p.`��A�`[Q����L�];�F��N�kITA�ʌ`�����,��wEt���F�r���AO-���úݰ*/��l�޸�t�"̐J�F���>G���gY9�J��6:\?�"7�־9����#�	�/���Q�]�xn�g���>��oY���ԯ�~��E��U���_;렱�|?4^�";c�8�+�*������}�7RYnh����X��IK�A�S�Zx�ߦ{�of�1Iz�q/?�������|��� ^q]�N5�� T�i���G��Z��a���&*_�v���%vkg�I�e�`�2#*uē̺s?�k�lқ���^�
���'c͹!	��6�Uj�����C���V�4��aF�9[�[c�d}P$��؝��f�r�2��D5�Y��� ��=�(�E���[�=ڗI��B��4������o��T�J�bKX4���(2�/W�D��g�1�!�K�|v�19U'���0gx.葳Ύ���Y�M0�^�Q���9�/���)�,yhC���Q�b`nN@��z	�L`����cJZ���ҝtᢤ�}l�S'pkBH�˭"h��ԿX��hط�X�c��j=���iٻf��9��4����H,�"�<u��/�^v$/L9#UN�(��Әn�=����(S���u�:��5[�[����ED,���u�(Z���=�w�?�u��o�QG�.����� ښOq�r��=?�\���oE�����6��\.|㬗оoiJ��qtKJ���n�����>��v-ը�7�ʭ��& 8"q�.�Yv;��޷�'�cv4.�R��F�|�$��=���c�k�tb�l;K�v�cWP�f��m�����<�q"�1ӳR�N�dh	�^��l+��"4Iu$���HJN��{�������9�������`b��kW��<c�����[D����O�D��x�qb�����~��/(��p\�"KF��
�#���0X^�y�h6�Dm��u��&�:��D)OF
�7�<>�W ǌT�%��b�c��Ѧ�Y�7q�r�y�MzG
����g�mS�	��[W�ɏ�6㡘k���h5mN��jᓘ����I�\̗���w�9��f�
kf�����,�)�XV���h.یm�c5��(cnb��J�����Ig����g5.�rdX#���ǔ��"�\�1^gC��ȠeZ�>�aSz���v�	W�v+)��d�=W�}{Hz�Ӎ���c�7�[�p������IC��.	��+�J��$��L�(���.�ܔ/�xF�ف5ԫ��@���vP9��O���&ECJ@-���Dhr�Rp1�ɵc�x�#axjv�1�U1Ty��H��3'��a�+ت��vi��n������[���i��K�[�)��ֻ6�������nu����c�5au��D�񨂘�i�r���h�ދ��a6��ž�[~؎=f%��R$���Y���ߠ�d�$��Z��/�ԆQ('	&�x�g9����H�N�t�w��-8���;i:LNFE�(��Q"���n<8�s7��=H���CMU�a�G�C�g��f��c��?j9\�ܦ[O��áɭ숢��b��}�y�Ѓ#�Yb��0v�M�?Y��<bAC��Äe��Xo�ߎ3�5�W�a�@�=,�����@ÍE-6��˨�����1�x�|@9V�-�R�������cK/�?m����P���������͎ ϊ��/[����Q���Ic�˾�@j�w]#�1�T�	�6"/�
���Lc��l֨��t�m�sTN!�,�T�B� ���Mb|w��'�߀+����4���ۿ�<||�~�`��^Q�$��eH����q"��W�OH�{lԐk�ڊs�'�Z��e���e]�u�1[Z3�����@���M����5ሽ��B����#��[A�ٻ�*�0����e����Ъ.-K8�_>�JK�y=��R����x�5!C+���Ҩ%�`��%ߛ��	�]�H�c�j��M�).�eD�TM�M�~�M��R��i6|�^���hͱ�Y�?���<V�,�)8̐<̛��'�u�~��7@��?��]��o֝b���g�J�^7�������rEy�y`	���E){�Q-��WM}e�w��/a�"XG=�c2@p �e�\p�I�K=�ot@�M��R����щ	����<A�dba�m5"ͪ��Ă��[l6!��gz������E�Jd�PŤ\�/�BO��l��!s��E�� ��X筀�-�K�Tk2K�'d�J�#k&���DdT)����#i|��U��<'M�-�Dm �pb�7��uBD��uӥ�����N�A
�f�|��1&C�B�@� )�g��m�@mQ�S<�'휭��pSH�(�'h{s>��w�uB��Aq�-�fX��L�Z����Ev��8;����1���ڷ����_ ���//��kq�"�����uf3Xj�k���n�վ7mv墳OZ����BtՐ��3P�C�r�p;:Q��9���N=� �G��ƪ�؂\�G$M����1�1[�[I��,��q�Ch���b�7K��/�Pr���=��u��3_�W��Mke�_xVpc(5J��T�����Hro<8�Gt�&Z\��a�Z��~��1��g�ϽH"=s���u��<�%�A_�xG>M��P�M���*"!�'�uL߈�	ջnL(p ���������E���:M�ɲëI1N%��� �� �����-sn��m���:�mCQgM�9����i���w�S'M�ۇtv��)kr�"iئ��A�_QW�����kB~�x�o�5�	��fs2WcS����3w��)&��1�Yc ֥�P~�MiRC�m��$�^��h�_8�f_��7=���S6f*/�M-�/�� g"ף��!���Go�G'*8�C��+�/�	��Y��{V\��|�� sXOB��W����R�g�=��Ы�8sV��������c4�����u�Rz|\�6۽1�K2:n�R�3@��5��J&m��d�{.�tc���aI�V��8��2Է���g����
���U�^��`=u��Q�#�(1�G�1w��xS�5��ڪu���x��@��\�(>8�I81�t�mm;������ւ�ߣWK1.���um�[��9��һ���LD.�j�b����C�"�{"���a�cJ�7�8�د�����a}�#�y�y��j���F��Tؗ���Vw���Ob���k�?�?�l�̵��-l�ya�h��q�$���ob�����zg�1X��K
�4�9������ï�͞.��|�O;(09K���5L]N/���E���R=�i�=����b�Dk�w�]���&ϙ���ޓܛ.ƺ;��6ke����)�M� �m#/ZZN�W�pc_��S`�'���C�<�"�q����6�N-%Ȱ���N�K(߇��Tt4���9ׅ#]"&�/�n����گr�)�me�aR�=��.4���>,|i$P<&��)�����T�py��[���o8�!ܾ��?����ݽ3J��B��}�G�!~Kk��M� kN*���y(؎b<�����8!a���'�>9��]
��k����s~���w�!.������t�������Tc~[F�j����L4�˾��� d�����	�m� v��z�Y�\�vb�<a��,�ka�o�m&+3�c'�G"��b�1��^�f'�����8�$�������DډO�Æ?3�������ٗ네bE��y��_P���<��(<��t������v���6�೨fШi�{��ӌ�8�	�,�����Z}<O�ko��r��4�w�+�L:vE�W�kmT��������v�ߐ�Y��3���>�xS5��]R]t ƺ�E�@�ߦ��ҭz��$	'8ѻ��?<�N=�^P%zG��L>���D��k���&!��sU9P���B���* ��IT��ي��$�F�+\�F�S�"YLaV�aR�MK��۶�k�!H�[R|��&
�ƶ�g
��CI-Hx,&��FM
ǂW^^���u+�ݾ_s�V[e��kbf
⁒��Q�ݳ���Q޻D�Ql]��x����k�I��$� �R��Ɉ��aj�?�ef(������>����j}IX�0�U{�^���[���wWy�������m�z���F/�_s#zh%喪|�i��<s�#zGd�P^����	!8�ι���n�q[Ά��Xe[;0����m�3�� ;Sm�j�N������y���iEQ���~?��U^�� �M�;�����f]й�l�鿾ȹ�2�
�9�h[�C��qQ̇(1EE��J4��}�����~A��f#�O2ң�L�Jz7q�P�i�ݪg���?�\ʮkt���7��1��,�m�أ�j_�>�F$o%�B��p-#�6+b0@��dTo�Gi�ܾ�Ʈ*5�X�I��z��=<ᕘ�Y�Rg��M��Ѭ���Z|��4�p�����9�L/�p�(	�����rit:�N�j���$c�-�ݱ�A���NLs.E�L#>z2���@�jHf��q�*\���52��p�\��e��N_G�X�s��O��N;lo����T�X�m'�/�{�EZ�&���"P��&�F���X|�8�z�U�K~a4j�C�o&ܗH`��6�W��KG�O�������H�B}�Ex|د ,�0h��g<�Yi1�lV�h��"P��&f��I��V4>/�J��x��E�d��ܘ?�ru28_>���+38�jw��Y9<\�cǌ�sab�eLL�ť���PH�9f�ڊv2e��v�ya�ʬ^Iy6���JC�e�1:t�7� m�`�����L^�8|*k8C��C~��_0��b���e�{%��	RQ��6���)"�3u��	���0�!XF�*�U��~�ޮ�~�G�H�j�%"8�k��ۨ��Y{���þ�h�cƍ�� ��\V���7���Y;���o��UUu�e���s�\W��m>;@��>�[��iO�q)��SG��gO>Iw.���YYqU"?v^�aXF�v,�I���ކ����N@�?m4��%ſGj���/n�M?��4l5p�͊�����o��-���EA�xw}�Z~n��e��7��'��5NSJV�ų���0��q��B��x`˭"��3����	�6���6S��LS�7�?�S�Ҽ+�.�9���OP�3z�e��u���</�����ϷTh�mɕc��I��QY��Ȼ�Oa�ޚ�;f�� �-<W��ˉ������#9���c��5��sST $�,�ѱ�S���e��'ZB�q�Ng��@��aZ^X��p����U#��_�2�Jc�Y��Ӣ�bM�t{��	}H"V��@�{4z!�(5���.�VDa��	�@@%2��|63��y�LE<\�ݣ�Z�Ce�۱*v�P�W4��V�jpSs�7_�u��[��p_J.�Z�3Q�q:�At�[��Th�c�pRL?��Y]��:I ǦDr=7֌�#g�ܰ�9B\���}`���Q�> ]�������fmZ�p��a`ptӤyڥF��4Ϥ�H%����5&V�?�<x�h�r��K55��1&�t�T<��\��SNC�� ��W�`~�e^7����7a�����R����fjI|�|@r����׎�h���4��k����1���-��a������N�_����"E��ێ��;g\�V7N���ﹻ(*1��,�V���)�а���ᔕ��E�@��O&I/�&,�o�d^�Ӟ�ܖǬ\hu �ǳ[�`Ù�l6) d �:��o� �z��c\�?<x$*s�[�T�Bg.|MԸ��������E Y)��(�b ��!2�>��`��q�gn��G�HA��K����eg߈%,N{�Ǿ���mNR��O��&�%�ts� ܧ�Ж� �&�����2H��>'ƙ�<�H���D�q�sF�9�9(p2�s�M>��Sm}���!�
�!��a��~LҰ��>i7%���v��ră`8����q��f6W��u�x���p���*aj?�˧�.�G	�գ���m�yTI�k�&R��\\��6��2��������Z���I���k5�ZΙ�`���cA�@J^素����P�q��H��Ѵ"��b5����#J�K#��-)�����Ug��r���̀�
x��*�gSw���쁘>�1=:c��;�bX(�>�1�=n�Q�ُ�!�\���p�j����*>����}��m��)�f����5b@[�B�U��o�~�Y�NA����ȌdMd����̓_�V�� ������ �w��Y%��$B��m���`�٪���Tio��Cژ,�u������:���]�וg驥��������^[�nm�G�'5<�H��N�G~�>�_3H^=�Q�v3_6rn^�WץI����� e_����yf���_.�G�`$\b�v0��l��$sn�`\�_5199A�}���i^p4$��B��bM� [*�K���C��ь?a��^�0	m	��V����ur}����zd�Fs<;W�����>��=k����k@�ɔ�U�.�$����>Ņ��N���ٮ�ߗ��`�6�
jo�/r�a�15���1� � >�S[.�'-��x����[��3sM&,<�����'�*�UcU�xP���nH.`�c�}t�V=�o���i��?t}���d���.e#�$a�-6٠�"��G�2�M�]V
�_<�����{؀��Nm*�{��3%3�)`^�p>������/]6
�ed���1�ɧ���a|�
?��(�՛���L�	�'�O���j�6�ǎ�LQ,���Ǣ����6���gReU܇�=}���ѧ^?N���}�����rx�\0sy+���Nm�n���2&Yt��f��[ݩ���47��ş��"lzߟܪ�4��0��[�_>��mj�lOƗ�ь�O���� �e0$F���kR�7����I���t�C���b��趶���A�(f�����Ľ��
qؓ��ŋ�@����ۆHB��s�Gv$h.���MR��5�%Q��`te�LzdrT�Ć']��sT�(U��%%�i.���i�.�G&
���� i��7�n�����`�����6hT�K�պ��r���V��:]�7��4�LY�֡�w���e3�Z��E�w������`�5�_���Z������7��9>��k6< �=k:ֻ�c7ޮ�4ݔ4�ZNTZzJzy���{Z���2v�T*��I�*�*����s����:
+o�s�xp�,�O��cR$¼��E�<R�������3_ -+�ov�(�6��zC��J�v߇~�y�����5�6��PC���p���D?ԡA{E۠��i(�=�_�܉�-�0�|����ߪ��mj��7}`��)��D�����m�����(\tM;�Ƕ�sn+�F��� ��G0��os������?D^�jWa�Giݴ߶������>̤Ӱ��ȣ"*^uE�]z����c�p>�a��prab��3{����'^A,�k����,�詰*!y���;�Ϋ恺Κ^<B}b'�|6��U򘂌��,�y��8 D�F�$H���e�,����ĆP�e]g9O侎����ǰ���lv�	T�b�'P��+b�EP�"���-^���7ƓY��U�.{4���}�g�:�b[�ϞE*���h�͡�ڞ[ߙ��M��_�w�[�/��_���V�ݵ�`�`:�c���{�D�h�at?��ӈ��Zq�ƕ<���Ǐ[_=��#um,6E?x��#�]��6���&����b>M��A'�v��G��c9p� u�Z�Wn�30g$|�{g���������]��=~�D� ��K_��aN A��X�d��L^67���tc�8\vbuv��:ocedpRO#p��FF��خc8� "�c���1�<�m�T�-h�'8�׵�gE����6����C)�5/�SKu�9�&�F�Xӯ�\�ׁ�$��k�1��w1R#0R;.P.'_�=��\�&>&E�ȑ|5b���M[u<�;��h��(�[ˈ�ܑY,&`�ڵb��?�w��Z��a�7Q�-��d������P.*����&hf�8��y�z��E�Crn��#͖%���U;"8+���c9q�w����F��s�͜�]8{X�>t)D��,�A�
�¡��0��j��/��ĔnM��u�@>��X ���fЀ�E������|�d]M[�&s�T/�]'�4���GE8���ϱ�,޵�q�)wϞ�(��^gɪ�<vm3�Cܿ��~B�����P1P '�/��Ջ\�@^�B�k�3�Wq+�^0fx�)��]¼s��\���	SH����u��^(���[�*��a�[���*�ǩϑ�G~�޶C��s�b�S6f�H�������},��:�=�Q$����~9~��q��q��q/�d�R0���;̭�gdU�R�Պq�`�zb�Q[��#!s�=�dގ+p��x�R6���ʺ�Q�}�}iK'tf$����ú�2n%���vB���:Ci���������9��]�_�6��<��g�1��x�k�fk��NEQ6���;�EJC���v���b���1�*��ϓs�D�c����ٳ��r#�9�yӖ����CQ�sؓ�� Z��n9�o�*̠��������t��]<.so�GF:��L{ �=\._U9�]���g���Ha����z�&#X�b��մ�뮨��6��q��H�M���냠2&Ɲ7��<�$�,1���
��o�py5���4˖��#��BP��-t`3��fȂ��˯�4���c�L>P�p������$�@��,�soQ�9�^��iJ�������@@\�a13���ˁ�b4����MY�V(KI�1��P᠊��lq�UD�]������1.�"6I/?R��?�W���$<]��s�1�����m}h��|�~�G�[/���oP� wv|������|�Ì~�r��Q2�a[�'�����%JUO��i��ۼ�4;��}�a�LJ��ʯ́��~Lh���-'�������漑�b�-[݉�j.Ū��]c��'�����G� y=}\�|�fύRk&�`����2�^�u�o�yt�����:P�
��\�����b�ԁ�Tr?�(G%d����2���L�ؾȠ}K�j��^K�IHdi�q:t@�����6�-̒=Ѳ9i}�f�b��rif�;T��j;���ϾoӴ�(�|�0R���VO��,����'N�G���ݜ������`y�_j�vԇ�������EͰ��Z�F���e�UgA��)�p1��H�n���˟)K\k$�N .u'����4p�`ˡzE��T>.��W)�ypa�O���y��^�KQ��\��8��P�-+�y��
I{�fN%�[6q��-��_���|��ޞ�2	?�1Y��BW��@�Xu`�Z�Q��$A��E�n���Y���/5c����gxt�ީ��G}�_��R�-/������<�V��r'5 "�ԛ�z��S7a3>�&��A���'�����F�W�;z�>M��pd9�{��f��1���Y���0-]'$@|��
I:�vv
NX9���E�P�*�Y���7 ��YH�\��"M-����p^��;4���3c#�Vb�� )U��JP.�z�@�Hɯ<氆�ڼ}��Wd���]�X�m�f��t�h,[Ns���/����"� �~�4&�畄-KE[b�c,<�� p{�p�f�sh����'t叄G�a��eN~@m��@�zb�ٝ����c��[��i9���7r���p�'<$ �� b��FЯ��"lh���Å<��w.r�������:[�Fst�N��F���4��<�⦝�|�[�܂y�qu�g^?�&��7ol�{^����R�.���{N�i�?gYi��@�+j=wp,u�l�Ќ)�5I�RGo�5,�->5����?(
0���t��|]"Jt��Ǥ��4r40���a�F}�9>p4�W�#B=C beJ��n�>��B(�
�'LSwI֞��9�"�
�w_����oji���>I?�*Y<���J���(�0r�F���ƞN;([6�B3/�" \�V5��� �bY+Y֏�]�6o��T�ދP%]
�2�@���:��9J�!�|�y��d/�������Ŷ��P���űm���g<_|�>�w#��;	�&��_�4�����5^VFy����xa�tE��1������9��Z�j��&��V�/-h�URV�m8�����������/�c|�2�V�~�����˪E�J-ak��H�A�遜8+e49P�5m����A�����kW9�a��w�*;T����H�zl�q�)�O!ٞ�!�|��<>�d�?.�M
��X3g��/��;����!]'����<{�÷hK>�0|�0^Y�-S�Ȯ_���Z��<E\��=)'�x��i����=!5ytI n�D��N�\���ޱ�K�'p���}�E�uߛ?hB�r�d�<�������;�ȇ��)Û�Z��?�|Fvt�Sj����UEģh�`O^Z���^o�"FV���np���qh�a,�5_���?� �.:^�u�ҧ�	��xʘ�"r���Fn[&k:�W��Jc�*�w����r����{�[�ˋ�������P'�6�tA�5�Q�����*��ȑ�n�ןe�o�w��/g�����o��âQ��u$���[��������r�; j�������W��m'g�p���$\��nx�qQ�����N���p�G�25)�sT(ܬ��1���>�Y#�HM�,E�IM;p�铿!B�������ʁ�� ��
3���!c�¡y�v �"��B�2!Wx�ZcP>�B�x6j=��
����C��o.?�����-Ǟpݜ�����`����5�FD�xeW�g@���:[�f�~Y*�}�/��<�9�9�D�IQ�]�V�������A��� z�z��B���"e�����|�^�G*�����J��B�;��e}�z�=t;ٝ�Ȩ����s��t�,qQ=�_Ǽ9��Y�)��v//Α�D5��Q��Q7މ7<�`����D�T�:h�R��oy(M��d�p
7�b�vC��W���ڋ�Y�f%�"d��3����?��~�M��H*��0��I����
��M��RA�f��������^��ۤv�;v8X�oA�����!Sw��Y�n�^��se}�~������2BwAtݺyO��+$D��aً�E3�w��l'\:ڹ�|��U4-���'VM�v��i����:�Dx���o�Χ���4ӷ�"��Bk�*}O�a��;hPR
���<�f���>��m5�[OV|�՚��}Ri���q��ї&�A�Q�y�o�Mܑ���4Y��!De�Jӿ%�4^����9Li)���(���P����6�l��T7J�T����Zl�+p�=�|IΆF� 2
D��,�Y�� ��)��d��_������m�g��q�uX�[
�f ���6�{�s���ش�8 �☉0��ާ���.�E��� 0�2��ZW�)�+�2�}�ˤD&�Թ�J:�5lP�����������o3<⍤i��u��򙪋� n��nN��&	D	�]�_�\�� ���2p�O=�����c*�t\���ZֿC���\
;�� ��6C_�x�X��h�XxV.���|�q9V�7!�(�.&���p�c���	Aq�͜�������N*�d��N@�B�d�uZ�2%���^N`��T��i$r7���
`�����-�Q6��7p�^��ލV5~�8����7<嗝b�u�s9��3������/2 <ѳ5��q�m�D�r�qQ����Qg���˸g2���m.��Ã	X�����7����O ZX�.�J�_t��TR�\!�RA��Z�"���J����,���.{���"/t|�k%�s�Cõ�U��X��s�rSl�Y
Ԛ91 va��U:���a �m׿^_���MŏTh?����%Z������t�ئBCSVA��;�*<aϤ��T��R�,!�= �a�y�Ws/���ƪ�����������΁7�ʅھN+�=���ARae���D�k$d^���G���*��h`1�~Y�a��w��7�Kh�&�r���U{���ӽ�WaSx�݁:/���s�k�$�e4;r��%�УZ�fJ3#EqL;�"��O_�9�8��&Dj1��d�f
�3�C1)f�>^9-_�R`��W�6�<�#g+t�8pm�C㺼R��j6���u�_�<$i� 8����b�ʷu-C��\th6&�{��q�˱����c����RK�it�V���ԁ�[��d���ŀ�^*VeQT�{�Sd��CJGl�A��u{���}�\�x�ϝ���L��.;?��=��q�,Rw��-Z��Y�>�_4�n�@�DFp�>v�9�Z�fW�M��:�5�󯱮�gn��l�&�h��)���l���NP���{��DK�4��;bi#&i�j�2�$�v��+�e��kB��.XR���t�ua�#��|������X`7���Z31�a��?浿�,�6t�s�a�ǡ�v����M{�Y|S���}\�*��J%֜�r���f
,�� ���[�H�������ə�,"�S)�{�g'-�#��6adO��߈V�ƙ�2��Y%"�U��е�>k�"�U��m]tl^t��/�n?LY��:R?���0p���B�0��)Y�,��p�q��a��P@J��'�!�X����JĎ_���ܿ�XYoJ,�Р�j���v�����` x�{�"&�o��z빐Yrxl�^KҘ��6"�_�<���\O�Jٜp�)Fĭn�	x��g����㳀��:���n=J�$k����Fl[��s7�`�7Zsx�eK��*��K�Xs�pJZ�Z�pN�q��U}EO/�K��R�l�JHzI�3��;N�u$;t�=^Kc ����@t��.�WH�w�����Vs��� �%���< 9�{s��gĥ��q�b[�-�Y*�T^f���ն$�w	�w���9�ؾrw�3������
D�σ�A/
�F$v+�=�=ߚ?�~�.pBq�P�͈��wU�/�9*��ajD�J� !Zq��;�k)���S�R�S,[*[�P��jP@0���W�vSq {�v�,�4���O�
�� ,y�QT\�p���pM�^�����8�Y}��=E�WjN���6d�F�l��F��_A��g�#YW�4����H:a:GW���+ő�'HaJ�� ��RR}!���.�v�5�4�YzhSc��{z3�oP��Ι�������*3��c=���0L���N���Q�o�ȶǕ��U�;���B�(
oN��<�M�?�v��u�*���ҥ�^�Amn���{��u��p�}t#/����S����	!�j���!c��_)�� �
�CH�7A��{�9�M���?�?�XP���#��$�gPĲ9_��ө8~��������!a�=g�D!:�^����[��w�!O�ة������)�HP%����Р�������g�+(K�7���������.9T1�jl�zH#�6���F�џ�]�3 Io�e�ͱj����6yS���p� �Ǎ�,�Ċ��K�X�Y!We�t��LW-��f�Q�p��w�G�72�}$Gn�hv&�,�;�I.�Z����t��= �ŷ����ʣB&ض��!���F'�ku��V4+��	N�dz7u��L��,1'9�8&�D��;��Tf�q��*?J�;b�MG��jl�t�ō��O�{J�w3�Hp-d�%'t��xrR�m%��we��������L���n�$��C���E�z��Mh<᪮zrv��r����H��#U��`*):�Z��^.I5r!2�@�$��FS�0<�� ƚ���w\�!���w!�.�l��}'߂�W)�!n(m�ѽ:�eܘ��J�A�`[�l"�Ep��1�o
P~YP�uM�>`��aN�T9z���#`a�eT����Y��H���C��h�Q�xgZ��!!B���p�m;����t�.�ҧ�.�kQ�iQ�i�9���i<�RT|�eE���}qZU=����I�Z2H�fp w8�P9�`���;l���T:�6^ �vw��P�>�cB�)�|�ph��ZR�
�$�e0�T�Rx��4�m�7�H]=���&<��5��э^�<~�)�/_,��#�@WLw��w뵤]� c���	m#���0=���j��<���)5M4��40� ce��Ot#�3��RCD���P(^���s4y �6CʗYB���&�|���fg�n�<ԡ@�#R���Ĥ��*Qt~�^�p"�n�?R��
��� @VZ�ӦDC�{�``a�!ĸ����ɻQ+�T8i�h9��>�k��H�-n߲�H���;���ߣ��0@D ��8��fߦ�@����tR�lx�P���4#[�HA��$ء�f	�2Ϋ��;d�=Ox�2������J�����!����`\�n��Tl�vxZYFL���T�@ܾ�U�&��W�%o{�5@W�ɘP�sU�ߗ>�l3qiIg��򟣿��b� �)D�4P� X�6X�"(+����Y��ܛ!���@]��m�]�Z=��ý�i�k�s'�C��'
C�G�4
��� �ĵ�>��w�bs�<H�5;��&�]8k$P-�X6�^9L��#x�G�L�Q���
�4�d�¨`�����"���>�������H�zqA��V��}�����١B�g�cŮ�㔰���a���������:n����A��#��J�@����m�=<G��Df{p�^ԟ�7��"�9\�������9QB� �����;�����!��F����I���?���~��E�zC���#k����ޓ����2����O+˨��s�J���U҅�����!�ts��2�0h� �$�
���VA�u�����S�H� RY�f�c���Z2D� �?MD�>S�Qf�٬���%��%�u����}Ѿy�y����&}���}�nV��p@�),0�� /풌L�H~1l67�o�\_I�s��k�\���Q�H�=.ĖB�6VR�58��]�X���!���K��l~2}	�.}�%=?�N��� �x���RD}�j�u���^V�HAԠ�T���-�X=�S
��5�Z�K��7!i~f��r�_~X;x������s �`<�� t'�N�;���b�Y����|�RԺ�
��m�4�p��XxO(��.).��	���%B��d�d!)��3md�(}���K��qw�a������G��%�M@Q���F������M�@�6�����r��t�`֧�r�^�4� ��������k0�z�n������ˬ�1��q�q�%0ީȼ%�G3����c�'�v4Rٯ�?w;*�@�W�z���/�@�Lx���'�\�����1�����u[3�H�����<��۳��M�q*}�RS����4 �%�`�ţ�蘕�P5�F�P�n#�l��pP�K��b��$,������^LH�O�C���� 	R&�"|v�������t�.d�'Z9i�	Ar��@���ҕ�
��J�X�(���DA�]��j"n]^ ��;:�_��%�42�� 攮oV$���*c������O����2{1��C�Y����P�f[�y�뮳y哟F_�yh�TB*o#�J�>o<w���7z>��&n���;��r��0�{3f�k�$�*?�>_�x'�?Q\[u�;���G�0QL�ض�)o+m�����@09͙G��W��;�����Bä"g�b|*�*�S�1q+~g$ �����`D�0|�vx�x Z+�:zq������Ε B�VU�lN�+IZ����°e����h�2h@����*� �'U*�tpae�p0�W ����4�
���5���Q��G6O�b�k����GX���+����D�zIv��d�|T�LZ_a�
����;�P�d�D�����~��Wr�)p���2�t��Wm�.�V"����֣F�P80}86rjJ�ִ�����9�
�t���S�?T�x��8��R������u�I�ܿ��9�ƍ؏`�Xp����>'1��rU��Ŀ�F�Z8��S �|�,5�RW�5=�{�����ݧ�����1��[�
�fbMl� N���N���Fu�%zMq?�Aфv�����f�T-
״��z���P��	��86��`��nHb�׸�ָ\u��n�\������,���S)��~�a΋�a�\��~�`��LB���3|ώY��0��c\-���;����ыv��8���/#� �
�XD�k���ų�?\��"*�X���GL�F匬`b�ߎ���1�ϗX��:R����S�|2�8��,�ه���Qo|���|S��{��ߦ�j9AmI{m��>�>�d��%�3K�
�<�"�l�z�_q5�bmyG ��Y���Ŭ#�I�'��Q�R�p(%Z{����Jz���C���T�S?�
��Rt����~nk�>�m��(Y4�
c7 �Hf�'PC{,�3(�c"�r{�xs���d9f�c��2�Ӣn&wm&�� 0�+����8��(َǨ���^�\z�~���Ҙ��Mn"B#¾/��m�V.7
��ܶ#ˊx�%�a�實��?)�Q%��*x��}��?i�kh�BU�ށ�d ����2�?�/^�n��q؃&��V��%0u�Oş���~�-k���Ț� �#%���V�U���F�
��y.����*�}3���Z}O^xhj����xEl�u�vR78!��	>�4��7�9v��6ϵ�A��Z����҆�Q�2P<���a�^QsЂ,^4ަ��+��6Jv
�.ǧ�w��r�<�d=���ma0@� ��«�Xa�K�~�Wߍd�<M����~?�膰����L�ځ��G��'L�qi-4r�E����E��U�� /f�A�
/��S�_���;A�@�1{*���0��>z2�\�WS��r�o
2�H�c�v�ɑ�`(���?�,�<�%�>���
|�'�B���������Z�R�Ly�!el=�6� ����p�B�d��>!��T!�����v�l��q��2�˺E_�e�C�ړ��i�YO0��Iq��D����#p�1�n�FS�/kh���eɕ�-���s�b�Q7w� �%~�;dp��#b WD-�	�����$�6���ҷB�k(5q�4 ��g�7Ŋ��IG�eL5�^�<�rb�R��������̙T�^�S��U��"�C�S�x��e"_,���Y�L��9�E�I��4���"~�^�xd��j�!�(5�F�ײ0�+�?W�h[$�8`,�߄]e�9|pAD*4�EѮa�Z�F�؄��q.���j�A�"W$��6C ��i���C��b��T�@��~"��c�rΞ<>�3�xd=��Y i��N�U�9��6����K�y92h��4�b+U�4.
s���D:	iI���(��Y�|Nb߯�17��}��F|��a�i������QZ T�)2����G	���9���]~7RTR��@|�1ִ��WJ�����I*��"ـ�V0�
���
�ph&_,�4n���G6@�#�;܈�v.FuQ�X
��M���6/�Xo�un8p�}����c"���ˎ��l#jY���e�
��J!�N���E�#�7a�6�'�S����&�X��}�*��J��l�/��OD��8M�� ������}������S$�ݹ�*�S� ��:S�d�t�*ƋL������,tM�R�@	����X���������Y�\F�!�}�T�n�o,g�"�o��0.��cVb�+#6�l[�N��0R0}2�e��ĶB�U�]v~�*3+� 7��b�޵4����_����B䭑�I����x<߸͆�x� ��H��H2�� ����7:�d�q��@�)���P:�j�":�c<�Z���xS�`��}n�6e�	nn*��1W��C)+�0�}�X'9������YIN
3e|���m����j @	���7Ͽ��4Y�r$�O��s��p��b��,rL���S��"�\(xq�$v�0ƾV�h=�"�ma_�CG���������X-�����eYQ�V����.��K�Y�` �/1����tQ����*�/��D���0��
ެ)���p� �%�+."�?,���������(� ���#�)H�twwwI��t�tw�Hw3�1t~�Z�O֚��g���;;����y�$| �4��R�v��������t��RBb� �lv�O����Bygu��c=J���̪$���a�2��Ύך�榞$b�F,��l@���H�5j��^F�����H�X7.�����'��'�3�L�b���F�_m��ss���H蓡�ZW�?c]�Q���?�	&]w�k�8ކUj��%~Wq��m�$e�bxKI�o>� %��O�_~��9��m,��6�����1d
n����́��Th�9^V	#3�ꎎ?�=���r�4-pc��E��]C���(�������}��E��wo'�~K���x���,�|m��ts|˘�NF[���ol���S�uw�4F�����]Ђ�0hΙ?�'�%��_�6f�_vS~I��_�*x׉��uBf)�l7��l��1��ޟK����g2���,�GP+n �Z~E��k��{/k4�w��6}W���i ٿ)@���{�B��ݵ�?`�h�S}���θޤ��AZ�A�z��T�x�͙��!�N�����qwJ�� ����i>3��wOg����j��3��s�B��Zj����#��:<����+8@t���jr�Dw����*w\�,��w�T�*�L��A�_���*��Q��� ��Jt����\y��oPX�G֊�)q��X~�_p}������k�ʺ�%:���F��t�5��@������ƒԋ��;w�'��J5�uOױ'���IԘ�3{�vP���q�5��E��Ӊ�a����.�A{��	#��^��H>;�N����6^>��wlA?��`�-���6C �ޥ)�c=��ƜS�S0#a�]~�k'�.��I<7ox�qs�����)5q���H�� >�yF+��hi�:C>d/����!��!�w4ݫ,�7��(�m�gdA�u�.��+� n�E^L��m�L���/�9:C\H���W���72s��� �)��z�Al��O�O��˂��)mzQq������I1�)8OsH�g�m��ʟ��u���A�{*k1��x=�����3ڛv��*;��]�PZ+Z8뫣Y�}�r�#2i��Ui~u&E�	�σ?[>V���M|B����ue��!n��V/z!<M9�M����l��>��v�]�3����^���F'��'c��:D�_�=��:o��5(��7�Ynb�ē�� �wj�W�o� �"�+3����68w�p֤2��C��)���{��'�x�Nc��̄)���}�CJɲ�9$<<���H"a��[�.�|	M�}����.D,��g�h�	�FZ��.�w8S�^P�ɺ�$y{��uP~Z�곗���z�{��2����D>K\����mFkD���+{?Ȏ{mO��t3���Ϭ@}vT��%`���u�{+kz���p/fCA$��Ϋ�0���;�_�V�]�)���#�Z�����[]7�v.�%V�pjn/6�0����Q���飼m�lN��/���;>~�3�����X��̮����b�����g�5���֚�{{l���Cx=�+�2X�r�v۠�����5*}�;�q1����=��	ݺ���
Gi�p���������~ty��tG���=�+� Oݜ����k0�(��=��{3�/�{P�z߆�)̆mhf�?����qf�u�hP8�s���cvĽ������3�����v�9�����\����O��������wϣ�b���Ы���r"Ȟ��:fUܻ28Ck�n�׽iG��rh#�Mi ��<T��,�{�AӬ��\�X�.S��Pm�A_x�wbx�}�����X��N����c)�>u��m��&�MM�(��I��u�ՍQ���H��~�}(�������i��^I��T �.��o&\��زRz9r�(0|ގ褧�1[B�XbM2j�l`��_uB*����lC�oO`��F�m���}2�_���PI\��*	52�枩���
i�l,B��~�@)�Ⱥ�@7���6;]s�J�,��T`�}���>�҆^��4VD\,�Qb+.�JMM�'������nC�~�w��x�҄�̂O
9,�XK���(����l��!�o�Z���6�����ȄA� ��\��o�oy��Ղ ������?|�@hU`C<�YC����&�V)I�E�C����&�1�XT��N�3�[��14:i�W��f����@UN�tz��E���
H0���7���'�t-t{H�F[Z�U��G+T$���y��(��?/=��P�8�C?K�.�(V��GX(y���v�YE����U���'�6�˲rt|=d7|��X"�L���B9X��i�H�:M�@���:���.���>��I+71`��R�'�F�U����I�[Zԃ8�
4F `��o��I�]� ��|qq��u�C�U-��=enAz�:c'�+��vY���\X�w�����ll�u�Bͅ|��S��e����>n)�N�+l:��*����￪h��Z��<a��j�����5�˪�Je��v������WPk�ÐWCTm?�t!~���/�?�1<O��2�P'B.ǎ�`����4ʻ0XLI���3�L��r^K�T�c��k&�"5^��P!m~�O��I�l��Y��Ym���t�&�Һ�I?F8X���c�����"�2�.ۼ�SՋ��e�aiiI���_]�=)�������l��R,�*��p�'T�:�����&��|䏅x)��O��ۭ�e\_4�w_��4NIi�]�����s�ōڅ|�/ݓY��[�=A`�?�Voҧ�C�ŎI|um��.�������RY�Y��m�F~)�0S12��P3�l|�"|�u�Cc��A6l�@m6\,+M��;�p�r��p�I��H��Λ�l���ɘ��+�$��q��R�L��?|/L�iD�D�vt��\�'����ol9:{�/��7�%�����}�%R1Ǐ<� 
5�C�V3P���2=�+a_�N��M���4�:a���n�P�8��'�c3����ر���C|��[�D-C-��4'8�ty�\��6}U5��X)D�I��_��7[��"��6݀j �#w��)R]��/�ķ����L����Lv�s��לk��sK�<��D9�c�����r��D��E�r�_��QZ����(���Ùp${���7�T��5�7К�}�'�x�����t��Ӊ����Vڪ1�.�@@�Ns'�E�礧�@'p�ٌFЖ�Et�	c���z:�G�)j��>�zxx�m2�~͜aB�g���ׇL=�(��0��P�o�u�[�8�~�Ե�/g�Ϸ$��� EK��7�zS�0���Hk�cJK�}�l��G+��� Ǐ���`���6�=�4��1ó�/��c�ɭ���O��}�N�' ��4blܐ�²뷱��R��"�"H��-פ �$e=-���+k�ӗ���Q:��A��jK;��j���N����6����}�9�Ӣ���/0ZgñLE����u�^�ƣ���,y"%t���n����h�6�g4	�4Q^y���'X�
WK�Q���'bVc#���_�G�5[�+%ô��0v-`�ف��H��Y�q�	�X�>���u<W�՗s�,=�����<~2�G���?�+����*�"������X�d���~/:dx~�d��-�����������fX��y���]�p;��UTI��Û�OX���e%�V�x�ԶX�<7�G�~�ͫ� j�%�B�N����4�c;uo��Q���o�;v�������5��Ǘ��Za;Ul�jd��"ە�7XL�[�������l��ٔ�l��]���ژ��A�i�m�2_n�4&��y�qy�����g�PߚT�02�U���}Pџ����+������X,�e'�N��g�U�Y@��&+S��lw~�V������I&�'ҏR�C��.���ݴ�A��Ѻ�"j�f�]Uo����랿o��.�o{������9 �^T����Dĸ�P�,�]Z���r�?�!,a�W�yS����J���V�J�������s�>�L$_n�fm�$�J����S�ݥ��5k"�Kt�uq�zqt�*` *7m37I�6G��9�Z
�wH1- ��� ��ES{�*������t~x��-NҮ��G�Иu'�\�-��/� �Ob2�w�SM��7a�P���,#w���+G��f���]ל�@D�틀ye��	�X�r�~NKSReo�\CE�Q�V��������w�]�jq$p��.N�k��v'�s�աoك-tt�iM?&�rl� ;��	�-�Pz���*�n��?�* DmG�n�+B}Τ���ar��F*�ѿ��_>P�f|�Z�SQ,:��1�L�[�7.J��U;��,R({�S�{U��y���d\a|��g���'LP�L��}r��W`E���\���o�����ܚ�I��.ٴ sa�y�g���rrdC�Pj�:����]鱗V���)G�P���A��i���9���v�Z��<���^�=���7�$���:s!Qg�n�� w�����Iq�N��m�*.�n�r��͆�)����{�/�OI���ZT���坡F���E���o��K�.�F�duGM|>|i�)�Q��7�����w��y$�~�o'|������Л��d'+EZ5�d��^7��U���!�����@���G�����\���baڊ(R��N�>�<���@����b1�
޸���а/ �w�V񭪴RD&� q�|;�-�=y�z�L��'���,�����7f�SzS��?��(�I��wn�Vx�F���?�C�O�j�i$%��W��Ν���� ���qcv�D�TeD�?�%���yʌ�V=Ln�n+�WMnQ+T��V�۪���j�")�f1d�9?��JO��<B;()�Nގg��C|;���&oAtN����n�s��ګ�Zr�M2��xo�§�����Ү����BC	AF�N+�+5'wwKyC$�f�MJG������XK�"�*&<��[��d�_���9��i���74�Am�;��rf���13́u���n���\YR�V�y��l�F�qr�`�ң�Չ�T�Ի�H�i��{���E�z��V��YU������"��~�"��DJj
~��2?Y6�"���(9�g�(�V����:��Ұ����1T���Ԩ�_���f���\4�� �2�g`q)w\%��5�S<��:�g����m�[����O"�G5�J��䲸�)�/<S'����J�]����KIS���[+�4�Q}.�gn=�
W�:�dҪʉ���D�ț�M:޷ H#F����d!�����}ܸ���>��`�d 1Cݭ/7��y~rE���fx�������w�)S��ez
�����z�����Ao��=��+��+��p�~���6�_D~Lx?}�fs1�? \�IO������H�8�sK�E!68b?��Li���𼌀-�G�b��BGX��t�Q-ĵ���������Jf� ��;�����>V���wK�X0C����TH�M*A�|�S]���cļ��?̆�l�\UI$��7Yi��e�>2����X�P<r�B�h�,���2F5n��0�0TT��UJ���w��
]�퇙E]���S��5�ld��_Jw���|p^5�)_��H��WC�'�hѷ|8���%|ѹd�>p&ӵ�����跈&1�$R(�5(��@�QH�jq��fٖ\vvD�h9��p!`�/��k��cX8a���5�-�.��H��Dt��=�/w��HT�[��8��@&)�oq}���u�W�y
�8�={��aӵ�{��lU�E�C@�m���/8��67�̶t����a/����bqJ�t��bP���{��%F��P�~��2����s|�n�>w'�~��F۷*q�c5Z�>��8.�'P�v/�y�
wT�,�N_d�g��0���&N.X�y����(H�	Z;ÿ\`���S<�E�n��z 4�i�'����Նwӈr�Z.Z̉��4�|����I�\I��C�u7��Y��CW�@-.םr��3��ٽ��m��y�]󒱨�.���t���
��ٚ�#Sie&�������c������ht��3R����r9�>�D�~r�J;��'���B�G�	;)	:�G�\m�.�d�����lW;X�3�o�о�(�"\ D+!���:���bZ��a�"\!__eS���8����0�A��{K�s�o�?ݎ[�X-Ӧ��bCt.@��O�U�qi̐Ά�LO�|v��g�w��/9�C��Wy7�u�*|(߱�e|K<MrQ��e��b��2wآ���yA�MZW�g�������;� ��,�P�Su��}s�ꪚAE���U�@@��{^s��S��
���0�
xX"�3�Pz{*�Wy��~���7�H���e��*�����lY@Q�]�%]��rN9A��m��2��o΄hW�5��1^r�>��#9#�'H��&���}�լ�UsB9L$\�1�5��n�g�\`a�J"2�n�o�&ZF�Z�p����tB.y��>�ݐ��@�����z,G%���0/ �P[KLӶ�H��R�CV�����e6f�q
m�Z��~�tpH[:�lf�!/�0	��� �x��a�<y��l$v��= KA1U�U;���"vi�nU��܊��0U'%��!y�q�C�j^,�B�T_KW���\76�o�F
�0v�H��O�ԗ���j���
JGl�˟�N;����PB���"��D��8o]6�
�ް#�)�l_����P��s�v�sh�1@�ٓ��.b:���Na�d�
����oxd&�eSُE�%*��n�+]K�H��I;5nW�(������ۖ0��h������&?�iH��u�Yp���,#��\n�L���� ��|=��Sdm���>ͮ0y"�@��K&�V�����'�W/<�����&�/��z�?�wg����F}�Ņh��N�_C��j�Ϳ7O�#��&��G+�q$B&[Ԣw�]7U>�=?��.?w��b����B�q����'�������,��ti�"���U�_z��
�¤�T>�@ϛ�}Z�.Wѿm��L�s
,&d���K���L�E��zհ���~詍�����@�^�Bl�ۇ��d�Z����/�è.�,9���Ade�©�e�(svo����P6a������ �F�@�����1W��"l��B��%/
�
���܁lO�Z�>h�$�Uy�h��-(�`M�m�sQ�}\����T	��,K�%Fg�R��]W����ƔM�+�6��v��y"����Ҹ�,T��u��tb���G&��}�HR���Rᶉ���Ȇ��G7���z�"Ϣ�
���7<4H�jz�y���A��߅k�9���}7�=Ts���v�+W���n��~m#��&�\k�L��-/�
���HQ�6`a���p�I<DNɈ(�hJ!��m�!��G�	[Q���_ku2g��@�e�T;����掬$L�Cc��b�԰�ޘ��P���q)3���h<v�U���D�dt��3�81<�i�'V:��,蝟�
�ǎ�����=f�/i���x�O��
��+by�=���U"ߦ�ު+�a�|	��=���fG�ܢ˫:A��7��WHx?����G���t�-iu~�%�:��3��6�#p�k���v�bl���xa��;{��Mݛf��@O�zT��u�O�Ñ!����B�(@ g6�˱�dzm��i����Ո��_���3{��[�0D��暥g��fn�#!s��n���&��.M�Lnl��6K���n"00ߎ�jx9�4�S9�RW9;���y����F��?w�7*F�E6�`��
d�5������K���q؛1P���;�V��K&��LD�|v?��e��4ɼ��_ht��%H�����fG��e�[TG�L��xݜBlEo���xd���	w�~�Z��/�����_�'E��^m�t�i�qx�	�����V��4}Ow�".>�B*���N����w�~w-I�_��e_�4�������im�%Y�!楠�?�����2�}�4��+��i\�ue&��,5�0T*)v(:�N�d�]��=�q�j�<$�@@Ⳉ�T�ÒC�ć(��.�|�R0 '����>��;��p	
(&��9�}�G�\ 9�D'�zWm6d͙���:��D��Ԣ�����3�"d��7���b�r3=6�������[4)��� �v�Kg����v��4�TJ�O�c�M�G�<b+��Ȅѕ��ǒ�qxZL^sO����vj/���I�aߦ�V�+���~^����B&+.�Q�dV�KݏY���j>��j��(y(4u{��Ut�4��a6[�N/�i��.ǲ���]�~sq�&��8(�΁4�me̗�&�6|�ۅ��~�����ϼ�BDW�ӧ��)�|��G�0���	��=pEiѳ�K�_�V�Sؑ��z��MV�.+�
fym,?[�k6�(��ܤç�㯮�&��6|./�T׼J��9Yt]to�R���mpR���{I��L�+J"�y9R�h���i���Q��l���#�L�9�Q��:��s��"�У�m�Q~f�	C8Q�����\�yC-*w���߭M��~Ԋ�����x���m��|�`t��3q�5u��U��j�u�¤��x����w�y^�x������}" �1��+5"�Q̿J�I�L�Eu�)b��\��p^��-�X��pkyp�Ov�-+϶Ȫ1��EӐd�y�Q�IwQy?[��'��	�,�Q�o��z�/v�_l���*�#o��g�v�����b�u��?rp3 g��F���QMS~�*FF�W�W�|v3|�\�&W`��TB-?y��v�uՍ����V�=,��[}�9�֨��I.�t>��2}׊{Ӛ�E� ���r�B�S3@T|��| �Ns�(R(_X`�z/V� ?( ᳴�o>ӈ���,��n��c�,y���+��O�������PZ�tG���o�`�೓�/�j�fzN��� ��<�]j2��vw�?�n �1�h��4���.��U�h�|ƚ�
/xѣ���a�
Q#Ã�'���__�>8��4��w��*�n��R,�:��/��%�]���5jJ k����v�Ř�[)D���Mb�:��է�4���S���wK� A�2C�ᙠ�j�a��w�I �\��a�@�ܡ����``j�S�����Ƚ^�?���V��yl��]>v����7��{�g�1�bH�aP�O�n�%0\��=�u�}���A�og= [���3��b��;�sr�דJ�YA*k;LY�R O4�a���dX>A���U6�3�V~���Y=��*�i����[���^��y���A���DV�rm^/3���afyt�P�w>��4�dR�F��=�	f�	j?5�a��O\�F%eh�ro�sH�욥uիʭ�tXgn�g<8	W�G\2WU�*a:�w6�B�Ŷ��vB�1ĩ��V^�.�u"�������|�ղ?���QKy�!��'ˁ��f�p<6�a������K<����d$Ý_����������x�P��gyX3k��?bC04��.>����9ڙ陽�}8�<N�L�ɩqL6�~����n(Aԇ�(@׮T�-P��n��}���w�=�hW��jPC�,���Chl)@�'�vU��;(_-`�dW��S\�����tc�=\%�I|f� >z�"��xۇ�wvD�?C��4:�m��>6�ߺ��r4O���U��[���kg��p-Hzj;�GTFz���^G,��x^}�Xڼ��z$Z��4"A����n��8��-���j1��5�X}�sk���wg�l�;~_���Kw�]����H��տ5(�8$�}`<͚Q>{�} �9�Í�~P�aTb����"�������B��s��d�0�R�s�:O���������y�Ւ����~6�w�aP��A3g���o5z�=w�L_�it�A��t�I����X�T��f��~���}+ ��X�f���Vk���|�J<d N���Z�F=�-��pk�p�;v(P�^m%l�E״���{{�S;4�<�^j���8o{eü��P���j������@<B^+g�f�k��!T�O*�$3~�kڲ�=k�=C�"\ŋ��!4�v�s�����f�fQo�~x�yVq��d{�V+��;������/?xc�Cŝ8w��n]fpkX��S��&�*����z5��>2��ۿ���0.�w�5n�����6X������������}�n'U����<�b�|��#�X�O�K���<�OʿW��S�1�
:}I;B�Js�K)4�:v��K	��x>���.��nh�����b�!�Nˡ�J*M*��'1�P��&�Qw�W[�d�J\��ʻ�R
�=C�DXF��e���B'	�s��
?��P�0�Ĕ��?�����xd��є���+�$k N�K�A�zT�N�wp�bio���*kl*�Y��op=v;��适�V|�bg�k@��Po��@�� l�����w��>�	9Y��|��S�6;ҜH]G�k��y�S�+ٝ泍s�
�8XKe>���n�����$K�k�g�Sc���&�aۺ��X��.�:��}fs0n�Kw>���l�(zd{��"\�H�ޘ�ӎ���uyT��*{{�K)y���蓈*�N��\U�-o��-^�8O�pbc�w��3���K��Y��}�u�Y�NQ��f�lv�=���7��5SJ�Ka�ru�v�7�t=��`��O1w��ZP��-+ I��q3�H�5��g�Dt��d��~�b�P���/q-"�E���9	ݙ"+VD�B��)t�P.��邿���&�Vb�Gu����e`���_e%8��L�=�x��ax_�T��� mJ�$�����v��gC�������������� �����j�Ϋ���W�#���O�"��0���X+{9*'������n�I%
�Nv��H�}���+5�)*�>����fgw����ٗ�OQ�QlzB���`� ����_uV��U-����; �j��"�D���p7���@>��>��^�~u�)(y	*����EĵC!�Ӷ߿�1��cG��^#�W����hɺ�亣20�l��bg�I��C�TVX���x��^�O�gJx�������γ@!:� ʀx�Lau��!����.=ʕ=@@�~�s��{������lW�	/t�lO{w��2bE�wa&�ђ�!V�ݹ�����:	`a���p�Ĳ�=�qI�CJϴ !���0��i��I��q#�qf���qƪ�5d9��ҧvŌ��!��N����P q�o�~�D��I�LО��{�M2�������/CK�̝њO�ǘ�\"�/ RtB%f�l�h�(0��M���;J�َD���F�ˑ0�����+*�%ĵ'�.���q �V� ����u�rv�X1�b�J~�oZ��$�挎:���� �r[�7�=�����C��*f\r���R�A&��^}:o#b����r�Yk%�y���:�X�l���5xxx�(���!] ����n�^�vL�|�iLڍ���'m��8);P	�a�����!r�4Ek!d>��V��4�l4:���s|��� ���Cw	�>�5�%[�%�����q�X'e~�����I�E+�+���}���7m�VRX��_s��X驙8��ͫhv���b%��9S
���vt���撷ݿ���X7�&�9J7i^�a4� :^�I(�䇟��N�%8��G檄�eИE�zX�� |�� i����%�Hulf�H�X��o����5p]\�l����q	g�x�+\�Y2�#��c�UЛ��_xP��
�;�#L�P�@��pL�Ƣ��i�X�k�q3Y��9C!	ty+�_��G5tޢ����*���7:("��������3RźY$�o[t燀Dx�ߧ�LH�>�r�ӭ,<ٞ���:�mI�1]@�B����Z�G]�hA��|x����B������_�"��݆"�B<�O>�>W"\�w�����ie�_&�f�ݭ�y��M҆��'�~Hc	f��~�v�+,��8��n�\�=�C����"�-7��.V,���TG����o�0�������z��c%�3i�>�����Izִ	���VҰ�����y+?���nx��	��2�w�?�H�Е][���4��1�Fg�>�+�ٻ�/G_ �x�8��~�T[�4Bő
)Ep�=V��Ŕ0N���g8�O���1fl,�>�`��4��bw�߳J�jXp��E��U�H�iRceHB��q��n�F]���1fPm�1����� F�"�w��}ֹ̮�����R;@��x8���K._�E�7�������U�M���+,�$�Ǝ�j��K���"��:��Ke�>��W0�x{'1[�����I%�KM%I�a�)ҵC�!����훥�L�8R�*�_�D�JIM���Bz� V� |�$��agѺ�v=~���yX鮌�������"O�]��}���I��<��0���W�H�䃻8z��ڞ�S7G���#D�졡��t�5U|��s�1e������t��G��f,x�l��׎Y�7�#w�+m�%]��aL���u����������2��n[vt��MX�͘�@!cH6�<����wkq�>��xo�W#vQA�",����6 j梘��X���vCd���	c-O��ˋ��+�I�zJ� � ���^�&����&�y�����
�+1���O���F1{�z���t\�K�/�V��
x+*|�x�t$��mk���G��	ģ#1O�����2�
�%��[�i2X IO������rĀ�E��_�j�wKa��:���w)��+�~�V����&Q5�q�)͟N�K������hy���f ��טq��LjS_�����?l�L��݄��	�ލ����Wo	B��c� �;��o9z��Aݨ|�c�
<)����q��`��0��D�|�ԙDsc<�jX�骂\mC��B��Iު���n�J�%��Ո�#�y�".O����jW��+�a�t"Xd�"i��T�ـp��P��/-��}��N��~�XB�2DC��Yɚj��L]I�v[9f��Z�Ԭ��^���)����&[Hd�d�]�G�r��_�]���.@q�$\�a���C�nH��O���V@CK���~��	��M7���|�o{rp�]	|h"�� �Yz�,@U�$!���Up�Aw ��S����$�KO(�h�����Iolr�c�<���L	����'h�g�����:�C��)��fu�ӈ������e��j߃t�pj+}�5Z-�%H��zU�R5�L*,ӡ*wζ�I�J�b>��r�yan4��KX��#;�Ǟ�Pr\�7V�,n��"���2F�h�r�w�{ER}��q\��Ws4�OF|��:�pU%q��&s�|�\��4ks�k?� ����~p��ǆ�]��5��ey��JT2hq�c���	���q�G��d�/yo]Ȁ�sS����������)�%����=48a�v�.L��«��,sc��#W��`��Ӂu�!���0��_f�<�}�u�n���0plgl�uq�B+�I�(�qbK}�K"��g1��Q� �Qf1*�Kn(�:�ٳ����)m��	���I1�����@х���L��{��7�~���u����xAn���U���3�K�A���ս>�3����6� ��cf�ݏ��Qx"�X&�y�z.qw`l4|�+m�l��z�z�z�4E�pw���ng�ux���#H#�pF�j�$pP�3�;�Hr��y�/�e,����'ː�'�Y�`i���_�����\ۧ����|���Ř��;d>W������\�ԾϢ"�>���t5��߲�p|��)����d�p��͜�X��ou<����:�a��}s���6hQ����d��%;?%��ZfZ��'N�asni��B!�{��|&8�����yW���e��4Z�2�ӷF�H,x���r�Jr>W}o@�� i�eU�}�H�*�(�$jE8�|���z.4Y����@[�|�]���FZX�ls��P҉�=�tq�~��:�a4�U�˄�T�'��,j���U%�|F��S�|{���;����]k�Yy����ͤ1��oF�r��~����`������Zl��q��ҧ��/���w���Dh9�^\����3�)͊�R�E�f�;��\�*E3�ƻ������E���j�N�,�ՠ����U��)��=�hqa_�q��ϝ��]���du�[RՍ�ƌ�ZPe�fpM9K�S�e|%�l;���q8�.��L���S�OvQ�,O�Rg֋�s4���{Ai�(��o=��w��	C��t.F��ws��b��&b����.bޕ���ͷ�	��ZF�3S6��	`���s��S��r�RZF�/�f���Ț.�vP��Q K%&K�:�&PZ��s�)��_Lg[ZԬ�O��9�^��I��u <��$��H*}�U�~�A����/�?�=T���2��+�/vWJN,z[�ǲ,K�k5ӹK`�a���
(�U,��~�Z2V�/z�53��|��%�����I*��Ԥ�|oD���Ru-���1��O6���n��QLZS���>�{�O�������VL�c�����x^�r���3R=ӸR�.�x_�W�b�o�-F�
�YxT=Z�ʱ����rz[�T��sdׅk�>�n���"�iZ}*ͽ���G�����2&�y��7F��م��U�B�附�J0h��XW)��֢3���S�2����J�&�H��WQ>�j�KHo=g�:��e�<��'���n^}�y�8@��:k��]���bi��0�\ٗ��s,٥�cx��3�W>�+�i�DV��>���8�2Q�p��+������eEK5�*��םc?oy�%�(�l�b��(9�*E[K��E���B�>�w���fm�>> o�>���)�Y�ˌ�&���U\�rK���ʼ����c5�V�H�s=�N���������y�b����8�˲ٵ�w��Ŵ�#S�{�5��*�`B��'IJ5� ��X %��q�V��{ky�n�[�I���\\Jb�`P���埍�D=-�^��Ā��*��z���Y Zѽ��T���C]n�Y%�d\�)1%X��3��,������,q�_�A����_�zrwN�.9��	h��v ��1������z�?p�PǍ���2�w�o�Q��#�_-1ȌE��EN��{��ݨ'4.֋���[D�0�&���\��I�at�Wx
�iI7D�%��X;=��ɸ?�ؓa�K��l������σ�+�u�O��z��d�
�.�$��.�g�1ث.6����z�V,Ġ�V��*=�#�  �O.���q�ȿ�������W��U��}��O�pE��l�~qF�Q�b6W��D v??^��g�#�_�Yz�4LĦb�� �Mj��`͆��평@@�*,��Y������,�䷖����	#Ũ���Zby2��.'�!�Ӽ���ӛ7!'���&��0�F_��v���6qP��9�c����S	N��8c��E��T�4�L���8A/R�OB���}��o�0��U����<�F(�<�#�0}l�F�=|�0�����MyQ P�Nu ���η�C*U�N.`%�욟ۉyw �-i��[7�8q*uC�����)=��&�� E��H�J���fZ]O�B�0{a��U��[مl�!~�9�;�Hۡ���Y<c�m�k�0o��G�f�ӫ��?�6w k���2���@b�5Q��JL2���!蟿�[#(�QZ��q��HЩo�ׇ0kj��:����_�Xy�9�w+`	�Rf24����GX��e+X�Ɖ���~ ���(Dqp�~X�ʇ"2X�|�%E�Pً��Z�i�X�2�ްrXlo�y�5�N����>�A��|
fe(�#�o��=xew�P�i�AU�$R�_����//�Z��f�\M帑�nsK3q}�Q��yW�"�VAn!�3��e4�RG|o�-ս�T�'�yx����̳��tC���9U��]`ykh�����|� r�Yenw��{;B����
�0""��4gm�L1wt�=8����@ q^��(7rY�?��z�TZwX������Rq��	s"*� J�"B�� ���t�j$}�sWw�sJ�Z/��ͧ�DZ��*����U���񁯴� ���GF����Kfͮ)��L%��D�ka�x�zX�E>;bmn P�*���[͋�.G����{�Ū~���2m���ZT�*�/��`_�?��e�%f�0��� �����X�qZU���A�Bl�Wp�wu���V��T���%�t��[9[���Nb�WV�Y𵁅7����¦d�E�O�}m>�]�IϚ�ؠw�rUwPKӖ��e���*��|8.S}xW#!�5�L�,˼տ1�9�10I?4��N�=�7!H~��?;'soր|����%^�T~d#�kWg~�� 0��,$�?��2��e�A�[p���Cpw'��{��!�������!��]�������#=����5������j���V��UW?��]���E�ԯl�C�JJ��e�����}	����4#}�I��1b �f�c1�LNĩ�6�q)_4��Q��5Q�"���60rf��Цu��g�Q��u?�L=��~��[�ji*�Wc�9]�>[�U /��-�&B�%�X�0N���-�n���jY�k��WJ�0@囅R�U(5��]1`3@�J���b��x�Br\;�>�S��ᖈ�殽Mz�qQ�K�\�fK�=�Hn�D|ګ��� ��������]W��P���z:�jl�ɥ�i/���N
��{�MB�ۺTh�?��E��M^"j���O�w=m:9�3��x�$O�߿	s�zr��:T���ǫ�����\K�#`�W�=v'Bkn���S���Ryw��6W�$�Ϧs{��!����.�J8�= 
>��(C�kQ�����o�������n{��JO򄹝6qń�o��b�%�gv糛�52�Rn�ǟ��5�cn�fir����\�,�Į.W8=sTΛ\K�;8�S����N��~�l�m1(��­�=��W�̣�y"�����ްy��i�!���X�r:z�1�s�+��V�N���:P��}�ZX�8o��\�+�	17O�+� �y�.��ҙ�Ӛ�
)s ��)��#���t�Y�y��5����f�/H#�2���\��[�S�t�^� @�Y=�jX�F�Wfs5ٱ�3�}w��VZ�Ja�{[3M��ە��s�O��+�6o�����з$Ɨ��"����Ő@�eM���{��o���ccd���jb$v�+��6v�%T�;�����DY��f?*��\�IÑok�Kz��E���Wm�8>I�l�#S�A�m��o�Ud��ʯD��@vN��|�`�iw�]��CRL�{��׌�B��/w6�ܚ,�!.3�<vVSr��@�->v~
�	x>qz��;�DvǇt72�>�f2
��$�����tg��XAy���rOb��T	�kO�!;�� @O
�]��� ���ro9?��ML�'�^%������V�*�l������j!g�vʾ��qqg�����A�B �w��.T�%�H���~t{L�:��:��	;"+F�������Jܿ�kn����4�]�	x�l��8���E���R�@ކ�MҎ}��tޣ��%����<�yOu�����;S���*�X�6��c�Z*��Ҩ��:y��ɭ����`�9��݊>���z�-���X��L;�Y!�š�� J<z�z�V.��=�Ԧ9�Z0hK�Ӄ^��=}I*�o�R-(R*Թys�Q��"̇lS��[}��d�`/�.�����8@�٧��n��yfY�h�%�6%�H�Y)��y�7�XtƅX��㬊m��)���߯_�[p?�O)�q���W�mO�)�E�:�
��.�{��j�.
����(Գ�Ħn�'�Gb&�/v��ୢ�}�6�Ǽ�"�P�*,��$e
0�����@S���m/��l� i7{��`j�W�4(�έ��D&�2�y�ˠF����#S9��
���%�/�gbm�6!;v�y�w�	-�)e�<��~�w˯�yEГWE�J�{t�N��p��-a���i��7��֦���O�13�Z��;n_(t�7���S�WJ��������x��,p9�_E��I�dP��<��Q+�������������fj�K2MP���B�s_g]��'v�7���z���Ϻ����C	��kb��s�~�[7�˾��X�Ķ���Y�Ht�����v%&7tq~�9�������Ga���/��|�L���0��u��1�O#L�]R]�,r��h���2��H�½�)}�K��d���4.%�������Ħ�y�v��������������*6�>���=�L"im��Ҽt�@$�e�G7����������f�l���J<'�+ץP��&q���N�iF0I��;.|o���7��3��7��_ϓ��<�.V�����Զ�-�z�w�I2G��ƈ�*�3�S����XaCO�>�(��fG$H���2�	��ǝ���K�Y�����/�yy�]�j��I3n�Y�gm�K�gd J�|I�W��3�p�t�Db��Lx��i�h���_T
v�3c��ʵ�}�I5H~?�ޡ�r�P�Mm���5�*>\��>4͈�[��v��	4)�&��\����`�;����d�NUٔ஻$*g"��ϵ4����v��i�C��Ш����zA��X�s�T�ZY�������?;w
�묨pc`�g���BQi���'�w��̘Dַy���b�)��6w3�,�����om��������"	��>ȜMf%�y&��H6Tj :�JFH��]��.������nr�勁��BXm���Ε�Ґ�����+���I��<Q��`,'���: �l�����[+G�m��Z���J���I#�w,T<�����S�G�L�j��NVJ�}�k���./Io��n�9�sQ�p2��NҷsW��I�?�O�0A�s�,z}�P�Ԗ	�L�Z�b��+�l��w�(�v��oT�ϡk��Մ^wh���0]�Y��*�ZMȕ��a.��gw����˿�.�dʨ�ߠܝ���c�]�B���Ŝ�8��a3t,kh�9_=P�L��6b��I&O*�6_2Ե�kW�99�χ{��O��)#g���PJ��6A��i�Y��/�lg'�\�w����.L�>��FM��HZF��Rx�*Ŝ�wVE��'q�/8�:��Mw2���K�"(A��p��ٶ�ol�S:�_Fԝ6�	>�we�Yk���;�D"Fw���ʼ�w�%>JN!����(�;�E�6�J9�s��7>��Jg�R!Ǩ;�B�B��k֊�[���+�;D[�-;ֺ�����Es��F�s��ࡃ8C�ζ
�.y����I>H�&k��sq�֓���INR����4�U�T����t@UO-��C{f�9����uz�^�EF�xg�xkj'��}0Q�.��6G����TDM$��Kp}]<��b�ؠ4�V�b��[�Y����<p�p�y�h����I���D�K%��`���
��.^L� ��'|:�6Xq9���k/�i�+L�]�;ʑ��)��u� ���qA�kW(������y���fE��TE�Ƒ@�lI�dZ� �	�>+:3g9���Z���ҝ�r1C�\$� �wp �G�5Q�<1�X�Xp�y�k��j�K.H��^&�Ȑ'_G�"��z,C��СlSZ�^�#�X�7��E��* �d�$ǖ����"���at!(ïu�������Zl3�6\Q�f��n�}w�5��5I����F��W �fV���3=o&�r����o�!�S��jѯ;|�5���`�'�嵇/%�_N�|ښ��/�h?4z��/��8����Y�%P�P��oO�Ȋ'j0�m���F�Gl�#�	��3��<��u����V�	�$یj�X#@d���X��L�<�|^ɮAڤ8���,e�e��|!o�0��Zej�|'�0�Q����@���-E0�a���3����:�I�)N�:��J�����6 �Wsi�jP�{� Ǟ8�ksLK���J�T��0_�ꍼ�O/p"p�TG�Fn���{lY߽�׉��&ڇ��cE����hW�o�2i�IzAÂ��c�z�2S��&"��	���a��i��y�7��gm�Z=�c�g��J��h�a%�|��kbJ�� ���B;���ڃ���N{��G���5i4��7��@l&(���1��5�{rj�����q�w�bVfSp���Ks� CJ�d��]͕�Y�Q3u�9.�e����8D@͛�}�oWh!'{�u�Q�(��Vn���J�h
Pw_���`���% ��Y���3���ډg2��G���D�6��	��[9����t��
j*�/'���w��8����!�֮���ӿߠ(d��v���4|��\�\���-Lm�g�H�u����R�OꚂ:�O��2�lV�w�
���C�I�����\�#�%:ۼn��z&8��Y���upCKO��
������L:b��F���P�A�@?a�p44�j����/7@�*:�S�p4��Xt�FJzJ\d���3�`��^>;���?<���d�ֳke:��ba���c*,9�"q*��g=��$�mc>b�a�
��	��G��=J�RkR�0�xX0u��0۠�����6�����'��"�)O�ACۯ�}���+��ϺCR~zΎ���/�F���Nj��Ȁ_�ʙ1%]���|$��i���)�9O�L9��?X�1�aEau�����HB>k#ݿ�����
��g�29����s�Quڤ1&wiYTG韷�f��)���b�J�_����}��iHtY� ~��&�z�y��x"�(J�}�WI�:K�1+�R�W߉٠_>s-��?��e���Sp���`���#)�j���0�2;�h����ih+��-��"J���$�<�F!�ǽ�O��~���ӊ���0����s<�aQ�ȝ�w!������m�� W���6o�w�D
�� s���0�x'�������� �o��LV�x[̙B"�'��x���&��&�@��}����@+�0��`��'�%�f��"��~���9��������M؟a	�I�����*'���M����Jب�I�^Y6�ݪ5c���w�(�GM_W��Y1�S��顕-�f���ԮMV5�J�
M����6e} ��`��_�cR���1��ڇ�Z��}%h�A!6��Y����>A	B��R\������,4�l8�4k{N��x�?�B~�����j����q1 ��% ��LK����Ђg�B��D	�h-7��jq�Ҷ;r���G�ɹ��̪,�����a1{xͿ�ڱU�z�*�/{�"z�Lٺyη0:���C�ڈ����`�����})=��z���硴���w�+c�~ n�Ն	�r1}gu'&|v_QG.�/n�I��`��/uX+��	��]%?&�g�+)�պ���E֍��������Oi5M��
	��z�O*�OZ�i�Y�����	�t��2���͡[^vu�a}�C��z~�m�͈"��@�t���y	$?C!E�bd} ����c1p�U^�٥qk���/�k��(�~ђ"�����aS1�N�&=eE�BI�(���=2=)Xi��7w,�=(�<�Dei���&�֡�i/���˽�hFydI�Uێ�_@q�6U���3;�cG7u�+Z��E����� ��̒3�����3B'\͏�����ӕᜯ*��'�x�M�0 Z�y&+��!g)�\㊦  D>C�bL'w\ b)���@LGi~9�>�8m���q��c�%{ݶ���BCc|��, ,�E�����Mua�{\�W����^BvW�X�X^.��E�81?��9wo�#*�ޕ��ݎ�Ǝ����ҥg�39s���,!��x���h�h}��h  �����'�o���w�v�Pect�(6%	�Xq���c��)�.VTT�3$7�E���ֱƌ+��nS��¡-%[�R�$��0��8@Q�󸒡��K���_�a��ӭ���M���x�a����a2�ѳ>�������|��ʮ��:Yb�s"�uoI.����FO�q4=ȐGbax�E+� �����b/Ɔ!oY�	�n
��Kt,�o��$�7A���;'&5�E�� �f%��%?�T�}���Z�9��z�f���E�e�Z�iy*�o���ԗ���70���˓�2 c�Ou�������Y;��E�gT�S��=�+]����u�דKW��B��!\LSP�aӓ;ٷO2ν(��p� ��-9��΀u��&|f�0$d��)�y�;�����-R�pgn�~!�=�܏ �;H���g�d)�q�ԟ���J�c��@(�����4�ɫzj��@N��1li��"��߰�h�I��ł�)�!�'�aZ���_疪w�1��#�|p��F`x�u"�+p���~�CR</=��"x�)�t�ÏZ�M�ݨ�5���1�qµ��d��B���(Mй�Ԕ{�F�
4H �!���\���s����C�E ?"��`ˡh�2��)��tL����n�C���P��G͋O�f�x��A {;ЯP�X��g"���U{m�O�/���a�.�3(5���7�^��L�5AM���5�m��v%��G�����61�ςF���Ur��"�	�>��^T�D��>���ՏIS��h��^��eh��/G�X�+q���a�N�X��*�䡊4~��*��h�{��T�E� ��t"�|/�!"� ^1��d�q�o�)�r~w�{t��	GrM�_����
�-r�����,R����_7/�4�l��X!�g�&Z�Uv����xw����v�W�`j��N�|G7��b�G��zϸ�KT V�<��O����0gM# `'�3l��A,��R�{`;�p#~֢��S7>�n)H l��K�(�KJ�)�ϭh���N9Ϙcu�[��^W�p�����5�Mz�dKm{�m8 �T�d:':���|��dA�2���!���dt#�[S�Q��
^8T�\�M����_(b?�$ ���_%����24�ɨ�D��o�����F�Ő���h��6��S4bۺ��@}g&Nԯ"������6��/ø� F����n��o} ��6(�#�"3H8?��)��>n����� �+@��N�U/	0Z��[����e��1#L�gIYh��_��Q����9��/�E��0k���j�P�@�����Yn���]�/}
�9*}X#}=r1��S}}���ڡz07��xai�ԮV�ú����a�f��v���ZW�����!H��T��y<��4B�1���uRWl6����Ko!�S��K��9�K!�mzD�-t,T�/�A�Wn����E[w��mX����~���=��z�0)%t�[�p�Ҏ�O����|��?ߜcݹ�%��������3��Z���mJcؙ�je���J�Ԑ�Q��~���i��*|�	���&��;����ב��a�0��U�W�\�C��:��a��HK%��u��̒�:�+?�P(�_�X�{"a��3�u��(���k��n-t��_�a�6T O����i6��Bi�g	�X8F P��$��'��{;0P�����<`�4�ڟD<���hcI>`��A�W�hX���A��@t��i���^�H0Xgg>(@	�pĲ����(cw"�����O�F/z�CSǛKX���4��Ӿ���
���:B�7��	��<���E꟫\��/�0el!�aGu��7����N�E��,�<�{�5[d��K��>F���F�&�a�҈���0 ��H��M�r�k�(_�(��q�ጦ4i*��Y��<dȆ���#�B�OA��r����2�v�H��{�Y�����3�Hl��t�~z��4!��Ƃ�J�ퟎ�,�,
�k%;������l;��C���t6(��o�	�f�8%&��@���ث��y��o:\��$�܊z�"�y���[��zd�X��&>	��(I� nL;��_����-��x�(ecq�eV���_yO%:��n.C��ɹe�O�k�U���]���DaF�?j�1���r'�+��#��+�oZ���-N���pU�۵��=6�#��!�!m�k5�٘z6��g��淵��|a���*I>n^��|!���ϰ��m�;���ml�o��R�Y�r����?��H�!��cb������iG�5��p����x��hQ~f^+��C�NA��3u�� �}s�0A��Q�1MC1B�;��Y�{�3��5�lMRݦ������o����gZk΍�ES�:l}&>��Ȟ3�����E
�"�T>��ϛ��ڷT�ջ���:ɞbbSŹ�Y�,)O:�g��6�W�
R&�W2�ak�h(�fl��
�h��D���6k]F)�X=��ʉ����V��s�Re��ڰ�i���I�շ�Mo�m8����nG��,v��h���ke�sXPr1l׬�<��� �H��i�T(��d׮S~�ő�"�S+��5fMd_�h3n#��Kg]m"%���?N�_��!��Y~�1]=�y��5��qbq{a�k����-���n0���o܅LT"��>�/�f��5�.���3��yB^��>9Я�of��B=���U���5ۙ�幮6�ڬxB{�S֮;�*�C�����0Rq��h�׺�q�qÖ����IF\|I��j~��;?�"�` %Ch�#4��El�-ӭ�b�uT�K�ݭ��.Xc��k/�j�2���XĘ�R{�1�w��_&�??=t��XSƨ��6+z��먱�q�2�
_�$�1�(�M��qP�$B�u_��F�M�����XTi����Ow]�f��n���@ h0������rSؿ?"�� �[d�S.Ƨ<�;4{6P,.�~�h��a(#��P �L����L�¶���|��.=j[�3�P���.�Y�ڭQߑ�t�ʬ���T<��5sY�:�"oQk���Q`�g���+�?;�g�ۢ?���s�D[D<��9fѿ�̴^��i�<�r95)�ؘr��3òl������������a
$/�[G��g���
7�.��	�	^4L�h�G�2}�\��wậ��f�<m·�ёl��A�� Mp?#�MZ�SRl��Hj��ު���Ac��E��'?�R�֬Z

��Tr���1��-�O�x��E���5���v�4�p\��i��+U�@0���b����mA�ދ��D�r6~���ǿ��oX��b�+����ϥ���Pt<sjv�Gp���иƝU������<��4�1�oHN�#�;��J��	��-���z��Ȣ�	�kD�v���������W�i�na수�#OZ��)��g�H���e�dڡ1�P�i�J��8��<�G����!���3���;:=j���v�e�R��ݡ����Js&�Ýv:�����%=��t�(e\����&0�Y�������/c�:���SA}QvB��>@�ڳh��CF��\R{r��~=����:d����sn� ��ܬpb�;T1����OɗW��(�h�8�!ލ�DaU��+���tv��I�|�&�Ϗ�?]BshM��7��:���<hg����_�?"`n`�a^_�C;�ضx�� �3a�l$4zPzů��NO̬�-!�D���S[�o�k� ;c�;>/�"T��݈��K���ɟ������5ncm��@|�<U���6O��I���419_�-.n�����i�DUN��@m2�%|�Bj-�� ��9���ej����������:�R�#8��a��w^�V΋0i��DkQd4�B>�4�v2��*��27�n�*�?����p�ܲY?J�����h��`�歁����JZ;v�����V�}6�Õ�z�����M@�nj�[��n�/2zd�T_,�����x���3M�x�ȕR}_����KO��fY/�?ˎ��4�ߴ0�Aý����*�A.�| �/�'Y�M<YRq�7t���*�������
�|�p����K,%�8Q��ў}�Ѣ:�y���%	��&����+N-��F����l�P�]Z��
��(��7b����-r���T�2q���0{X��y�>����؊>���r0���ojWlO�'���1�9�����QED�c��$�IO�Bu��oV�?|��;������PT;����Ny�B��׋�$��)�7��i�1ֳ}�)B�����L:��7޽�2��1��@�0휯�?����<$��X���\rw|�+D������҆xN};(����!�"UX�������]�����=(Y��`�����G�E� ���Xuv��-�\�(�K~�����q�(d��y�\�q�M
��^K��0�%5�ȬW���(U�G��=��&����^�� M��m�D���a�߇a��*4�Q�x=�N�Zr4.�2?����7�ޞ���\���M��Ȇ�[�aD�٫�?`3�5�zB��D���k�om�ǋEt^P��~�9�PP~������Wm�X�>3�0���@�ղw��&��R'H|A�H�V���kS�Wo����zs'�*�^��Lg'��R �D;U��R���w�8??Y��8���
>�u6�RRsc�x����m�T�ѧI�f6b±�t�B� �z�W��i�")���ɜc�]�f-�6�s@I��Ǽ�e�mIc����[J

�|�F�y��I�l�.ХxP����EZ���;�sv^tro���)8G}f��E���2�O|8��ˤ��v��:\����}�����&y�͈��Y�	~k��>=��F/p��i�%�D f�X���s_}��:˔�,�d�wr���=��b���O� / ;rȴ�0X�֌��֦ŏ$��&��X慸�_?�'t�^&�Zs�f�����<b����8�\�-�f5�Wl2q��2(H��O
�o$ X�Ӽ\��q־�\�_U�pI0���x��6j�5$e>�����^���5���?Ԙ�3�a��{⛡��]SC��]�·�5����x�=�)l�P����ie�����zHOx�gAo��) ��������
u�IQ�L1U�9:
�
�^$Y�4�9�Y�h���6}�&��z��?�*��˴�8�F  �[��bX�hx ә�[���A5]`�ޚO�lc>��/ӱQ�^',�u��-���q�����,g��WTd����s�щvjҬ�7��}��O�|4So���a~�B��H�.�C\�q��~��d�+W]�tb�T�����@�Yn@�Oڟ���s|rK�a���;��37��<<��%s�������ҝ�[h�*�������j]��b�ІA�Zt����͛�m�2Cc�(Ȣ�=�Թ��KFY��3`�Hy�a8������'�xV��K���(Wڄ�jϐ�P�����1.~T��>VR,č(�kw"�,#��Q(�syqq�}qbo��4�l����V��Q5�TB6n��U�GΡ�P��
�ٓ��9$(�:s����Z��:*|#U�@.�uZ	��H�[��rz�{G�7��
u��\�jQ7k
?>fu� ��������TX���7�n7�@n�U�V�I�LN����?͛������BV�ȡ��HCй4��I�	�J��j[%��M�0���4l��c>��F4	wڢ�[/�(�J�jX�����q_]�j7�d[r��U=�I�Vl0�v�ݱ�?����`�d�"���ps	�N]U�j\/Z)�D �̹��>�"�DD�fP��A���$�-]��no�e�Hlüx |mr�a4�[ů1%wA���v�g�e�Ph�[S,��6r%�������R5��ͫUS_&ú�.K]�J8D�,ϕ=�U�g�)%A#���"L���QK�%ݸ_�V�i���0B`D������(�K+�w�9�����R�n�뇄�^n�-@�	�)�:��Vo���������Q�#u��cr��\����>�F��=����Y#&;����Z�	��pZ߁�	 HԹ+B�����C7#g:�h���}���=��k4�=�CdrX��K���3 پ�*�˞E7��#7��2[�/��&�|��O��O)=�\ˆ�O]�nn�*��u�����ΝLY9*�8�hޥB�7��fn"�V�h����y���	o��-4���s�H�t��[�څ��7w9�A�W=}�%_��E��w���g�z��Д~�Bb���#7��j-�_��q����n�Ǳ[?1ϊRP7
NM`z��٭)h�_�Ǔ2�"��}�n��a�n��;wa��-�3/���+%�w����b��u�}sC�����5xd3�V�\�Q��-��m��n�J������}%Ole&���lr�7��7��樔!� ʤ���.E�`�WԦ��^aθsUMl�=?(�װ,6�	J�%���<�B���?�WE>��<��lhl&�?���X�
o�[UUR
r�_�jnb�:���ݳO�<�����kN]��)��4��Cp_ݐ������:F�z��?tG�jh���s�>=�d
��T_�w^�}�>�FnċS��'�y:h��ӛm��z:���|0@$��&�M�ǛVUΜ5i���>y*��=��Vn�03�?OJ袭U�G����4s�!|� *b���l[o��W�H���7���: {Ұx RTA������6槽�iO��}u�/�d<o�rU�<̊my+�_�bn5��"㑷o`Tbl�81�mDP�L�8Ě��l��Ⲕ�4�[Y��>�{#�rj�'��0-A92�#;8S��<H�9�]��.�'_�H]���!XG3L��	S���L?/:�[(h[l��70�=����z��|�U�)��.*��%E���]}���e�h_(��3P)<���tQ/�_&$�����JR O��Cn�Ֆ�lyԙ�C�/S�hQ ���Æ��T{��f2ʑ<��!�t���vh>1$����v���ڦ2�v/sh��P������+��p[4/�=I�u�*_k]��V�o5��P�6eӤ�O�)<�oe	=��T��g�HY6���~?k��ӂ�Py��vy�uSV��[�q��&��Tef�֞����%5�	���P>���ITL�#T'?*E�~��m�B�w����}P��gơ�����C���N# ��m �"�?�8�F�}s1���s[�7ɿ��@i��ζ�N}�z��3�
�X_�7Nn���R9��W>l�u	s�bw�yQY��0��.��Y���'��t��q��Sw�!���-��m�����9ɔ1����B���><�TI`4�_���Cj� �P�Ej���`�v.��#<�u�VX�b�N�C<���K��O�}ұ��TL~�ͺ��÷&�gTB�ҥ�ߩq���u`D����6sIhQ/0��ʢJ�+��i.@r4��T�"���>�f�8���<���f�~���CM��߶�����vX˖�p���|ro�{x��O��ӏ�J��/,����S�@+�-`�R�޶��%+�՟�&� \zLYϫȻ�� ���z:�Y�l��� 
�����[En~ԋXH�Ħj�u'�6��e E𜠍~���&���O�β�Q�֚S�簢�(D�����y���Gx�VFNR�e/$�]����7Ν�>��?ˡ�b>~�6��b��D��(VY����rbj�WY��k3<�Jx�&���A��V^]����\�Z�i=.+W����'��"<QV[�^�	��+?$������ 㷀���b��'T(���'�Ķ�_��?��<���S�����I�8�p:�vR�Vɀ��fYF6��v��E�^B6����Vc�:J�BKS@;����c.�g��1H�4N�մ��.��ծa�P�E�%0��>9f'����x���l��;��hl�?�~G����7Ff�!({��1��}}Uȏ�P��� I~6���C�b�hR�Y���|���0$�$]��Դ�ٳF��ɖv���Ru�,�|}i��[./�SΤXe����c�6�U�a����<Z8�B�ƍV����;���c�_l;���06����[�>+C�]�I��=��iQye/�ĳA�A������o:`d�D�P}n��m_�vA�T�]��S&ͣl���"}�S��
ܰ�&e_���f�bO�t~�:V=���R;[]�8���U<�T(fԛ����*2GS�}�(/��ƎY`���}�;>\c�N�տ�yL7�<��p.�?��ʞ�������m^�+�!Ku����j�r!~�wVou���xL+�![𧫁Ƨ'�~�K3��A�O2H��C�u�r�k��ݥ��F�术���|�.sI���й9���7�G���qo)W��%�`��9���>�8��Z��Į�$�|}c�۾��`��ܿ���<��~X�������7�0w���g,�A�˙s�iİ6_Ο�{*�Y'���:�Ms^��_���+�^t���{i¼�9#����L�xj����b�k��*� &���Y����6��CCCF�{T�~r]���2��&���W�⫠φP�Q����J��E>��ݢ3�<7��L޽E���~iD�J&���s�/�������a������=��
S�M�G<bل��2��ئI�R�l�>s�#M*�N=�!����4oLI�Rh$(Ԥ��֨�߶O��4�������[������k"J���L*�IH�������E<��(��锇��z�Gf{��o�B'���eԧ%������lX+e�ח� ����/3 �1e%��p}����}�t��Y��y�Zl�}���%/G�2�m�ww}2�ii��"@�c�l�b&��8"��խ�^�/��Ʌ��`!�V��@��R�}�剆�ୱ�����5~@ՃG���X��zB/�2���K���)ء�2�d5'��x4�c`t�ڳ��B�����ů���]jN����l�\�
���.�?x	�5p��Tݥ 2������&SEf�ϛ�����������v�&�/���<]��\Z��ީ{���ֵ7tP3�&���� s���A�8��r��y_(~^{jk$�[��*sM��=J (���av/fy ����kO")ISj`��B��8��z��o�x�^�dVQ�­�z��h�� �ꗂh�]��{�h�%��t��9q}���?d�7(#ԇY6���|���}@��.�`��Ҝ�+Dt��Ռ`�1?"<�mj���r�8^~k�jb�"�*��}NW�߳�Ak��i��c1u6����s?1�^�-;�ia�畋�nݷ>��k��*�Ŕ����	&�&�)��m8���0�="�4���αd�C���C�E�
�RRQ��	=���<.-��"��f�9�����(��#����a;hj`�o+�<�ѵl܉$��Exs7T��j��ק#[�C�����B��Ȉ�3 �b����hLl˖�7�ͭ3����[�z�A�>��P��A��М��m��],�z�������������u��4��8���D�JQ��x}?4�>���k�H�T�H�_ǫ�V�^���؃��<v�t���͚>��!:`^s۴�k\F!��o�y��t&$��Vt�����^=�@uD���F�&�1��1�Ԓu�D@��ohq�{�q��P�W�8�I�=B,��"��{IӘ�b�
̀��sth(*%���Z;��S�1�oY+�OK�<-A'���O����j�x�����]/<����� �fh���Ee�ʏ"�����1k�w���p�D��@�b?�_ b�l_]����	�>��;U�29S:y�.s��:��zX���6�Y�eU���
�*'e������ň�����:�^u�:m*I1Sz�5cwԛ+Y?6'�9�(�EՍ�
�'�o�Xڝ[} ���`��p�2I.\lK�5�A�0�n���My7;�x�3���8���MI�h�$*�Xx'���0�U�E���4����ז��:�<}~e�}0xէ���%�=y˸b���^�d�7)��9�N8��������=C��=a�7@�v��2	�-���s@u3�70��GgS�v����z���@W�ҿ���
�2�YJu-Ayj�LT�����gִ�k-��@�%��g�>Z�qf� dt������k���t��J[^�"�&�:@8�c����7zjx�������+V'�[hLY17}%��nV����\`c�=[��7�)��x(H�8
�>GAų���F���j��AG]������N�9��9��Y��c�j����xJ��^P�n�MC��'KK	E[�8O�9it_iP��\?4�^�A5G��#�_����{*;��x(�57��3?[~��p<�f�2��|u��D_�颭TS�K/��]��S
��̑��;�)���lQ2a��~;h2n�Y\�T�_����7u�|cQ�	2���\�7b.x����/[�Ҁ��*8�_�y�9�P���{�V����c�ޯ?簀�#?��`�R���D�Ìޅt}�1���3�ߔ:�B���,o_?f�t�ڋ���.�F �V��ݣ�)�S?"��U>�+�oJ�#�O��0��.��,�wڊ��u���`���5�߹*�0yX�,�.-N��%�Ƽ������J�A�_�[�w�.���>��BAQӰ�t�������J��@6нZ�pr]�*�nX���yZ~m����G��F����س[�\J$��a�9>�#�`�)M�s~�����#,������o�=�ⶊ��ۘ�X2��op�sG"	EF�;�qz��rK%�⸗��a��"�d�\bky~GȒ��ÅSvw�U6��8��Q �E]��eAy�.�f��ք{��f����xi�/,���!��V�,!�.�t���:��6�*V�Hb�rߜ�S��+:_լƚ:�2��v9�imJG,�$����*� �Q�u'Y�����{M�W��ߡ������M��F�=ж�P���3n�ۤ��v�'�ӭ����>1 
�V��kx?ğ�����+�[�`$��e-�� ��M��
���HִޓD����W�d�]��n|���(���}u�x37�H��ZZZ��Ү�'�}![��q<P����~�q����e)>����Ħ��~���#L']���U��Ç���U������t:�aw�A�~8�U,�K������������PD�J�P�����N��I)	���B�%����`��=s����/_��f��{�u]�^kOQ׸��O�҂�,��I'�>�pR#ϕ������]�I��k"R�(���*ϑ���W�i����&��]��5U2e0�t����co�����;o�cպW|���#��Z!�_/Wa|>�[�X9�}��pYX����z|'t�ӄ��;�6�ٯ2������C�C�\F-���U�z���t�������	�2��{�m�^P��K�m��L����m����N&ǅ9 �梮����Z�I�)�#tx�̸� 8��;Jn�]��-�FX��6�q��2�iۥ�gf�a-%Y��^5z���*6|(�y��@���
,�������l��o�N�������n"�޵w�;�4v�߅��ku�9B�����m����޿a7����K��۵�gR�M��$�����
�m�Z-��]I��&�̏�ҡw��v�0=��4�I޷Õ�P�"覃�*�������l̤^��C��~��<N���b�;g�
E:��.\�y	��;\S����'~�d&%�dg$$G}�|:	K}��U'b<�k��I��mZ��W��
��m/Ե�*�|�[-�.���X?<�Zr�ԉy�g���������'�0"buI�͟K��b}�j,��0��Ph�,֖?"�^���������٨qoh����e�����z&�B�ߊ�#]�<-h����A*/��������Ii�����Ir�2m8ΐ�^�g����"����M~I��6��H�j����"�����V:�!�NF(���.��4�g����r�������+b	�:����`*ڸu}w-�u���? ��rK�U)Z�އW��U2��U3w��"+/�f�	\d����Jp���9�+�����L���R�StÈ��~��@Eb�l8�.Ht��߫��7�K�#�5�ɛ^�R�N1�B�����*<2'���3r
���H��5f�zL�	��t�;�k,(�w��<��S�ݛYx��+3蝞�|,8���vǆMLLLU�R�3���:X4@� zCy�Q|��x$�&#�(�:,�C�XCDI�wH�$�ff4g;^:��Q�S�B]�;WU�Fȹ�~8۪JJK���:D��)��׍��� Ϋ��K7 �|�ւ�lL������
1CH3�nm�g�� Z�'{���ힹ
⓾��^��8��Ǆ���k��4�� V�l2�@f�@�y	I	qx
����+�m��S��=��fb�n�/���x/��v�	������o/S%|��^#��7r`�X5��k}oZ���ەl�}밭i.dX��xR�E�g|����fY[u�}��!\u�qq��(�F�e���`u��qR3�]mp��(�/����M��Q��Zj��%_���i�Ηo�[�?zR�#�������%S�2�m[��_] .6�]�C���������*������[	��k�)���I��D@@Ւ���C��t�p��.�/�/).����T�� t�5D�vf����O�{���e3�fS��J�;��R+[y��%��:�dR72�{C�OWre��"^~�y-�2i�"^����k����$�AvG������&�
o���Ӈ�ZLn��^t�}�/��|��f�aW�F���?�oU	�.]X1�\ˣz�lɫ�v�2����)ߣA��h�3 L�i.f�kK`��j l������`[��!�d�u����3[lH���EW:��}=��%ȯq�(�?�g�U��`gozL��\�EZ� ��%#3��qq<�Weg�LL�ω�E��8����1E�r���.Z�]�	>�� �ؑ^��Ď{b�l���-&��7M�X��a�}l�f�R##�Pr�S��TM��]s.C��%LJfB��1gs,�E����LE�~M�3��.U��(�>54��n��з4����R���u�}����Yl��T�#��������g%���#�1�����d�I|n�܁�?�h�p�5�j;���.�h�7q�&�JzVgFFbg˾9����Y6�)5J�b����^����0QR[oc'KODi������OT�{����VR�<E0�����g�~�%J�x1�!�����rZa���~	"{�VF�45d4Ab�g��'	=u��ݽ�c�l�~>�Z�Wκ'����)�:;�7�L=J�|���R���Xg�e��]]���{�N��v^�%�zUJ�H� ���Q�w�"�y�7{w���;H�.�W�'��=D�������v��鐋���`���PP۽��?��c��O	�hE�j[�|e�Սg.c�<����*@��x�S��:!<W/� 9"��<�ιD���H�`��}k�zh �{�|A����͏�ﶡZ���J�����`±���3�8TV*�L9%#C
o΋}p�'��oN�`�(�u�����m��z�G�wF��6�+��y����J�����}�6�d�	�6���l���F�� A�i�쑚��ao;�B�s
�n��""�̼ U��xlMԴI�@+��8@���y"n�����z<9�4".�񝨈�p�3��~��YG��ָSz��d�>"LJ�$X�|!��$�P0k� ��g��C}ڏ�@�U6���y*#�o� �3Ԯ�MZ<��<wR9��e��%��&(���j�I������>}Ї!B��T@���;r�HQ� 2�K�4��C�\�_��Zd��Ej��^�mƦ����7��-��|�c��`��V�i�M����B?�r7R^��0�މP��M��K2;n>ے,:e�~�:LZs?��_�M�$���{"疏
t
�j�f�������	��qu��GF��)����?��>����F��2Ui� � 5_����yE͗z����� Ȝڸ�+����'��Y��mX8�	ȏ��3�!�c���G��j�2��'<OʡXlЌĜK����̴\�r:ǑS岯P�7S���KK�u���^`�m۝>����� �9�a�Y�uYr�������AOh�Go`\m^1�y�1�[��j��H�l6�Ug���Bl=Ja�4&�����f^���r0���1�%%�40x+���Y0�W�_��П���c)�}���'��,��ƚy~����7K-���4�|�{!�u�	M.b!�%!��F~b�H?U�{\�"������m"$edB�E��4���G���<�)<j[��x��i@[@�6}x��8X�(E�6ӲL��낐��͇�4�:@��-RS��A�2����]}oNY�x��$߯��n#�]*ܕ-A�B	���6�ˮ���>#���S���/�N����8���U<c��?(�Z�oM�7F�GƹSf��g��f6�R �Ȱ&0�� |��\�ǝ�y��ͅw`�3�DƂ��;�)�3T���?Z�ѫε:�p6����3�p��hAQ�����>�_��21��w)�?�X���N���{�;~��3��P�f
�B�1XO��Id��n�i��)�i�����58͵��, �j�*t{���m1{A����9��|i�/��rzY�أ��=��k�6�2/*��˕��^!-�w_a���6�#wW���]��� �����
ᜯ������.wx/��<Ż�u��i��ϋ�pM�`�U�#�z4>�^��490tV �H&LHL���y��o�eT���B0�iVT�[CQ��'V�u���-O#yDȋW��Wх��B�x�2z (�Oo�V�6�?���|�0Zd{�]~7�is�  �s"(�/��z��Z�h��7A��o��� �rB�Z+m�&�����ߎ�^Żˤ��u>�X�v1�D�oؠ����,���E~62e;��ì3;��.�,�k;��`ZɁН!	�y ���]qv ���.g����5�c��+W�R�O��0t���Ӱƃ*������Oe{hr>ʊ���-^Y�5�����J��Z��}�u��P޺�ZJ���N����A����7ؒ]��%M}b���Tu[M`���D���V�e�X�Ӹ�x/�)���s�f�u�V���˔�w_�s4�'`z	���ckc�v`�.暿��j��[�{ە�<&$�
���AdwL;�tGw��`'�^ʊ��<��/���u�B�(w�L����M�&j��dj���v>�7-c*i'��pO��egZq	B�����62���ŇY�ΰL�(�e��K����[�&Iqx]
c�F0%�ț ��X~�b�"׋�U�a~���X���x�'��^"����{>%���4 nAKy�) |0���5�n�c]�М��Y����ֺ!b��{�m�Q�/}J��#��m!�|ݟp��y�=c�#1m�I)�?��n�����r)�2>��-���w�k�/���=w2�d˨�����uS�����@�Q�U����b�Vp:�zp����^VX,�h�r�xTㅐ��~��P��WNug~N �đ�<'E�C{���o�%�w�K���:��7�rH-�4XV��F�����49�^+f�Ln��Tx�������ab�Ψ��ه���SV ����>W�;��8e�g�0��e�E�Q���WRH>8ht��	�b3���}���g��O�o%�l�Gا��L�O�Y1�W��V�#R�/��U�˱�+E�CJNuz>ƎKį<�^��te4��}TKk	��� [��˘z��dGү���s_`N}ًD�;-�3J��-UU_�k��o����R4���-';����,�W�jc窄wb
}VK�I�J� M�/z�*�H�䂖
-���A)j5�H,~����O��h?��[�[ ����$Z�V��Nf����4��Sfv�e��8�-�S�1{���Ib���=[x;?$�fZ"���̙Jơc=���ɨ��i�Ѱ����r���U�����î������´��^�������ߥ�*��~TP��6�|�H/�zF�LTk�����=ȷ�-�ZYn+�cqb���J��q�䏻�����;u� IBMVG�l���*M�J��Ċ�"hsC�2b���.�T�(��|$LJRfA�J]�ׄ�_V��� �[�Sj@oU�b�9����ӧʂ�*̳u�I�D�5����("3�{�����=�1���Pi��|�i����dɉ�
l����%�	�R�A�*=3s�i�L4R�Wi�^�IQE�F�V^M������Z��5#�e���q��g<Bs{��܋ˮ�o�eޏ+��VW�W�>�ݥ?�k��߷���"��l��8�o�u|9f�3�M6$Y�*��QA7ݶCw��0uE��ֳ Q�3�6����C�&{w�E"����؃����y�L����UY�>.�����v�
�"T����`�m,C�%�4��AX�`@"��{R+�)���i�W�1g4�j1�_3�1@���J?�����'���G��l����M�w9����um.gݔc�D��w�h�5e��4D��5�x����H�+��7�Wb� �Q�f?�z�֚0�5�}jں�������9t�m�c�ζs���L~�[�$^E4����	�lL�K�d����{�V7XФt�4�����"�bΤ�����Z�ʥ����^�g�fl��=s��*_�l�߯����D���!%A1ؕ_�Ɍ�n��`�_�ǯ{B�_�Ní�{�C_N��q ��^�{����v-� ����l��꠼�uG<��	%7�� N`'	7p��&�C/��J"�;@%�W#oZ�_��O���юU�͚I}8FS��{�[Mk�P>��{~��uzPr��m[o�n�H�wH��!c:����~K;��AZ���TѴ"ޏQA�E5S������a�էu���i�5��]D�dS�El�b6�%\º,����)Vu��@,s붖_� ��J���O�$#���W!�H�:�Q�f�{�l61��:#e���i�L���x�¨*�w%�}Z��xl<�ɾj	��1�R�
#�ں��;<�"� <F�V���d�O��V6���U4��C$IeG.(�D��I�]�Q��?u�L�D���2J��w�tyKV
YflؗE?�M|�#s�ސÛ0�y+ѯ@Qx��ҋ��3�kO��>d�@ъ���?��~�U�i�O�{9��f�X��Ղ.��<��h�cĘ�:�| �"��xFR��N����� f���(����pbT�����Ҩ�+��9�Cu�R�[�gbj�˦�G`Glw2��ot�'��&s�֞��Ҙ����1Yi@Td*����$J	՜�)�MD�p���HI��պ�df� ��E%>�S<�ϗͼ[�˰� �eRl���;<�� ^~X*9;eNE=������7n8��o����H�Fϗ�	������A����z׆���lHN�1�������R��r�8}?/�N3����u�ݰ����r�Ʋ�g���+����;�J������׉�Mx���ð��+0��!�l��qsp�oX��+"�|�/rC>�Edn'�F�������6t���?fk1��}����9[�H�e[ۅ9`qThx8��;Y�}W� �&���w�Ղ�	�?�V쪴h��Gx��匊*����QXT2ELy5W��69�R�])�_�9�H�z<��551s�0T�X��������s�	d�����)%to���+b:Z��&[������\a|��gEx֨�����|R���s�%�_տ�`��<������+q�4u���Bf�[i:��NX�efW�vm-�=w�xC+��H|8B�5�iL ۆ��[5��>P\�#0(�$�|���Y���8)�vWfX�Z{9u%����ږ�����UF��w��l�����~v;�}E��]a?�Z����cP��#V#}��]�h�i�\��5�kcN���A�0�Jv���h�`��2���@�PL�}�����RsocM`H ��שː���O�g���X.y���
b�B�=�Z//�Q��'�٫�UP�)T������gQ"�}Et�=��!a}SJ��x�%�a�)F��L��J[G�����h�T2?��
�#^s'{��6�$�S�[���Pz���&�y�K���I��-��[`L��틁�~�	9Lg>����21-�.8��cj������������lB7kKP���\aJ���Y�	־m���_{��o��R���yq�a[JwC�`��b�����Q�GL Ď�gY	�$(B���s
��8̆�(�?��NH�):{y�
�x������d��-E�&�S���G�̩d���v��oa����"���dv�w
�l8��\��\�� ]�;:�A���y��Ұ������g��n���$�v���xk�W0} ��/�uE���
+4Eoy��KT��b�zO��s�ލ3�ڳ���CŢ�>m6FC�6���d�ؾ��	�Վ�FmEm��Sc����
B*�A��Uw��W�wET�9����۶R�! {�7�vG̦0c��%?���^����ɟ���^x�%�߿THo��f<`���ᵺ�8�������ھ��V����/vph���f�(sJ�h������r�r�1I�[&����R2��Q���֑6B��ȟ'[Y��sK�^>��>?��D��WF�yh��WU&M..�� \fd�:�	�p�����s������I:N�0�~��%�28#�z�O�/٣�)X�47�Ccw���v� ��cސ3s<Sެ�����Db�%g�.e9@B��u�Wc% ��ս檆s	V_����gb,���%���F��*��2~˯��ooM��rNx�٩cJ�[E)�*]����g�~?��yʝ`�\w�+G��o�l�/8�e%��
Ӆ�"�x��ڐK;����j ����|�C�q7E������]L�%L`�ow�9��/_c˅�=f����Jq�hun����8]��OlM�L�뽹��$��$X��V�4N�╢��S��53,�x�g���)��X��~��v0&���9�2��t�pi}�'0�C1qVVF�b���_�Rb֏d��5�iY��z�喛��1�8��=o������җ��I͸��Ғ[uE0f?K7I���#��R6�����d��������`N~Q��;�7�¾�G�\f$�s��s���R���'��8�;�U�����/���9����ƭ�[����f1�}��W?ό:T��Wޑ�ɰ,-{/�9���7����J�ʼ&�'"�b��C~1h}�X�> �%0���ۊ��Q�y�(W[�AC�ݩEv�I���vث��o�7%����g���n�O����Y</�?�
�MG��7jQ�z��GM�~���A���	���������V��S���1��
���s�rVA����f�JZ,�z�x�������D�����&A��.���: ��-��BE�5y�̔�9�q=9��6�6�o��EE���5N�\U�jo�˱r��t����Fqx�l�$��OZ��3H�oU������jz%;M�;k�5���u��l֩�����tXQ��!�_5mx|�.av�Z���0�s2���&��;���=�ɭ��k߀�1b����b��}��~�D�²�Ϟ�<�se������Ax`Uq�p�x�b㹇�a��J9*p�������b�K߳�|c���+"F�'�� ���"Rxk�e#�D��(9Z�3�_>�v�3̢�>-�<~��LCyN�Bo�h���h6m<0BW&o7oX�%¨��m�@�'L�>=z�)5M���ߪ���=�Q��|;�U�(X�o���{S�^(�w�%�K$���]Z@�����1>�m�t���|%p����i�j��1�KS��o/*�ɯ���9,-�x����7�;�8�Z�e��	��i�K�9�n/�<�%ޮ7-�n���~����8�ᬪ�RyQ�?�����mT� W@XVRXA ^�@,п$�=[	�����o��+�N���>�'����O�w�����*�?
���b@BL���nO![X�_�����F��Ҟ��G��￀6�W��7]�fcSPZ!�>̭��[�
)���PK   �kjX#���  1	     jsons/user_defined.json��N�0�_��:�|��;Dш#4ìFrm,;c'����M)%L7�hv�9��.���΀)�	��,�3�	�z�"��K95�����综˵g�&���UJS�77>�R�����s^ �S�axi��%A̔gM)�ĥ�U��Z�, �ٕN�0�g3U�]�����Ҫ�xع�T�Yw�L��w3�V�N}�Z�A��)�%�����c�l	�y���w���&|\N��f��M/�f5�j
�0X7�e��'N����w��rar���vU}�^�6���7pL�N�W���P:�G?x2x���G+}�?���w�6�ߤ��;z��l��O:�~��K٫��YkT�6c�I�5V��B��b�*��R	d"xQt�?��G��C�>�=�A�`Oʟ�ab,x��=�����Wy\�q���*�PK
   �kjX��vr�  ų                   cirkitFile.jsonPK
   ZjjX|�<�d� �� /               images/3718d1cd-d7a7-459c-8466-c70e7021b870.pngPK
   2acX�#�(~ I� /             �� images/e51fe3aa-205e-4659-a3a1-ad304791dd1d.pngPK
   �kjX#���  1	               :z jsons/user_defined.jsonPK      <  %|   